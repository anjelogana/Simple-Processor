-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Aug 6 2023 18:36:21

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "simpleprocessor_top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of simpleprocessor_top
entity simpleprocessor_top is
port (
    o_Segment2_F : out std_logic;
    o_Segment1_D : out std_logic;
    o_LED_1 : out std_logic;
    o_Segment2_A : out std_logic;
    o_Segment1_E : out std_logic;
    o_Segment2_D : out std_logic;
    o_Segment1_F : out std_logic;
    o_Segment1_B : out std_logic;
    o_LED_3 : out std_logic;
    i_Switch_4 : in std_logic;
    i_Clk : in std_logic;
    o_Segment2_G : out std_logic;
    o_Segment2_C : out std_logic;
    o_Segment1_G : out std_logic;
    o_Segment1_C : out std_logic;
    o_LED_2 : out std_logic;
    i_Switch_1 : in std_logic;
    o_Segment2_B : out std_logic;
    i_Switch_2 : in std_logic;
    o_Segment2_E : out std_logic;
    o_Segment1_A : out std_logic;
    o_LED_4 : out std_logic;
    i_Switch_3 : in std_logic);
end simpleprocessor_top;

-- Architecture of simpleprocessor_top
-- View name is \INTERFACE\
architecture \INTERFACE\ of simpleprocessor_top is

signal \N__7470\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7431\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7350\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6705\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6567\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6537\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6258\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5686\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5673\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5364\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4456\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4360\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4071\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3993\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3970\ : std_logic;
signal \N__3963\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3879\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3772\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3751\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3741\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3738\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3702\ : std_logic;
signal \N__3699\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3663\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3660\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3618\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3612\ : std_logic;
signal \N__3609\ : std_logic;
signal \N__3606\ : std_logic;
signal \N__3603\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3594\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3582\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3573\ : std_logic;
signal \N__3570\ : std_logic;
signal \N__3567\ : std_logic;
signal \N__3566\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3542\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3522\ : std_logic;
signal \N__3521\ : std_logic;
signal \N__3518\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3514\ : std_logic;
signal \N__3511\ : std_logic;
signal \N__3508\ : std_logic;
signal \N__3501\ : std_logic;
signal \N__3498\ : std_logic;
signal \N__3495\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3487\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3473\ : std_logic;
signal \N__3472\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3456\ : std_logic;
signal \N__3447\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3435\ : std_logic;
signal \N__3432\ : std_logic;
signal \N__3429\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3414\ : std_logic;
signal \N__3411\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3401\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3392\ : std_logic;
signal \N__3391\ : std_logic;
signal \N__3388\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3372\ : std_logic;
signal \N__3369\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3354\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3350\ : std_logic;
signal \N__3349\ : std_logic;
signal \N__3346\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3330\ : std_logic;
signal \N__3327\ : std_logic;
signal \N__3324\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3322\ : std_logic;
signal \N__3319\ : std_logic;
signal \N__3316\ : std_logic;
signal \N__3313\ : std_logic;
signal \N__3306\ : std_logic;
signal \N__3303\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3301\ : std_logic;
signal \N__3298\ : std_logic;
signal \N__3295\ : std_logic;
signal \N__3292\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3282\ : std_logic;
signal \N__3281\ : std_logic;
signal \N__3278\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3274\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3264\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3260\ : std_logic;
signal \N__3259\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3251\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3237\ : std_logic;
signal \N__3234\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3228\ : std_logic;
signal \N__3225\ : std_logic;
signal \N__3222\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3217\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3207\ : std_logic;
signal \N__3206\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3200\ : std_logic;
signal \N__3195\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3185\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3174\ : std_logic;
signal \N__3173\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3169\ : std_logic;
signal \N__3166\ : std_logic;
signal \N__3163\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3153\ : std_logic;
signal \N__3150\ : std_logic;
signal \N__3147\ : std_logic;
signal \N__3146\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3129\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3123\ : std_logic;
signal \N__3120\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3114\ : std_logic;
signal \N__3111\ : std_logic;
signal \N__3108\ : std_logic;
signal \N__3105\ : std_logic;
signal \N__3102\ : std_logic;
signal \N__3099\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3090\ : std_logic;
signal \N__3087\ : std_logic;
signal \N__3084\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3078\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3072\ : std_logic;
signal \N__3069\ : std_logic;
signal \N__3066\ : std_logic;
signal \N__3063\ : std_logic;
signal \N__3060\ : std_logic;
signal \N__3057\ : std_logic;
signal \N__3054\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3041\ : std_logic;
signal \N__3038\ : std_logic;
signal \N__3033\ : std_logic;
signal \N__3030\ : std_logic;
signal \N__3027\ : std_logic;
signal \N__3024\ : std_logic;
signal \N__3021\ : std_logic;
signal \N__3018\ : std_logic;
signal \N__3015\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3013\ : std_logic;
signal \N__3012\ : std_logic;
signal \N__3009\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2997\ : std_logic;
signal \N__2994\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2988\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2982\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \Instance1.un1_r_Count_10lt11_0_cascade_\ : std_logic;
signal \Instance1.un1_r_Count_10lto11_1\ : std_logic;
signal \Instance1.un1_r_Count_10lt17_cascade_\ : std_logic;
signal \Instance1.r_Count12_i\ : std_logic;
signal \Instance1.un1_r_Count_10lto17_1\ : std_logic;
signal \r_SwitchZ0Z_1\ : std_logic;
signal \Instance1.r_Count13_8_0\ : std_logic;
signal \Instance1.r_Count13_4_cascade_\ : std_logic;
signal \Instance1.r_Count13_7\ : std_logic;
signal \Instance1.r_Count13_10\ : std_logic;
signal \i_Switch_1_c\ : std_logic;
signal \Instance1.r_Count13_12\ : std_logic;
signal \Instance1.r_Count13_13_cascade_\ : std_logic;
signal \w_Switch_1\ : std_logic;
signal \sevsegl_RNO_0Z0Z_2_cascade_\ : std_logic;
signal \sevsegl_RNO_1Z0Z_2\ : std_logic;
signal \r_HexEncode_i_0_6\ : std_logic;
signal \r_HexEncode_i_1\ : std_logic;
signal \r_HexEncode_i_0_5\ : std_logic;
signal \SUM_2\ : std_logic;
signal \SUM_2_cascade_\ : std_logic;
signal \r_HexEncode_i_0_0\ : std_logic;
signal \r_HexEncode_i_0_1\ : std_logic;
signal \r_HexEncode_i_6\ : std_logic;
signal \Instance1.r_CountZ0Z_1\ : std_logic;
signal \bfn_2_9_0_\ : std_logic;
signal \Instance1.r_CountZ0Z_2\ : std_logic;
signal \Instance1.r_Count_2_cry_1\ : std_logic;
signal \Instance1.r_CountZ0Z_3\ : std_logic;
signal \Instance1.r_Count_2_cry_2\ : std_logic;
signal \Instance1.r_CountZ0Z_4\ : std_logic;
signal \Instance1.r_Count_2_cry_3\ : std_logic;
signal \Instance1.r_CountZ0Z_5\ : std_logic;
signal \Instance1.r_Count_2_cry_4\ : std_logic;
signal \Instance1.r_CountZ0Z_6\ : std_logic;
signal \Instance1.r_Count_2_cry_5\ : std_logic;
signal \Instance1.r_CountZ0Z_7\ : std_logic;
signal \Instance1.r_Count_2_cry_6\ : std_logic;
signal \Instance1.r_CountZ0Z_8\ : std_logic;
signal \Instance1.r_Count_2_cry_7\ : std_logic;
signal \Instance1.r_Count_2_cry_8\ : std_logic;
signal \Instance1.r_CountZ0Z_9\ : std_logic;
signal \bfn_2_10_0_\ : std_logic;
signal \Instance1.r_CountZ0Z_10\ : std_logic;
signal \Instance1.r_Count_2_cry_9\ : std_logic;
signal \Instance1.r_CountZ0Z_11\ : std_logic;
signal \Instance1.r_Count_2_cry_10\ : std_logic;
signal \Instance1.r_CountZ0Z_12\ : std_logic;
signal \Instance1.r_Count_2_cry_11\ : std_logic;
signal \Instance1.r_CountZ0Z_13\ : std_logic;
signal \Instance1.r_Count_2_cry_12\ : std_logic;
signal \Instance1.r_CountZ0Z_14\ : std_logic;
signal \Instance1.r_Count_2_cry_13\ : std_logic;
signal \Instance1.r_CountZ0Z_15\ : std_logic;
signal \Instance1.r_Count_2_cry_14\ : std_logic;
signal \Instance1.r_CountZ0Z_16\ : std_logic;
signal \Instance1.r_Count_2_cry_15\ : std_logic;
signal \Instance1.r_Count_2_cry_16\ : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal \Instance1.r_CountZ0Z_17\ : std_logic;
signal \Instance1.r_CountZ0Z_0\ : std_logic;
signal \Instance1.r_Count12_i_g\ : std_logic;
signal left_1 : std_logic;
signal right_1 : std_logic;
signal \sevsegl_RNO_1Z0Z_3\ : std_logic;
signal \sevsegr_RNO_1Z0Z_1\ : std_logic;
signal \sevsegr_RNO_1Z0Z_2\ : std_logic;
signal \sevsegr_RNO_0Z0Z_3\ : std_logic;
signal \sevsegl_RNO_1Z0Z_1\ : std_logic;
signal sevsegr_7_ns_1_0 : std_logic;
signal sevsegl_7_ns_1_0 : std_logic;
signal \r_Switch_2_RNIK7AZ0Z11\ : std_logic;
signal un1_click17_0 : std_logic;
signal \r_HexEncode_i_4\ : std_logic;
signal \r_HexEncode_i_0\ : std_logic;
signal \r_HexEncode_i_2\ : std_logic;
signal \r_HexEncode_i_3\ : std_logic;
signal \sevsegrZ0Z_0\ : std_logic;
signal \sevsegrZ0Z_2\ : std_logic;
signal \sevsegrZ0Z_1\ : std_logic;
signal \sevsegrZ0Z_3\ : std_logic;
signal \r_HexEncode_i_5\ : std_logic;
signal \SUM_3_cascade_\ : std_logic;
signal \r_Count11\ : std_logic;
signal \r_Count11_cascade_\ : std_logic;
signal \alogicunit.N_95_1_cascade_\ : std_logic;
signal right_0 : std_logic;
signal right_3 : std_logic;
signal \SUM_3\ : std_logic;
signal \sevsegr_RNO_1Z0Z_3\ : std_logic;
signal right_2 : std_logic;
signal \bfn_4_12_0_\ : std_logic;
signal \alogicunit.un1_a_1_cry_1_THRU_CO\ : std_logic;
signal \alogicunit.un1_a_1_cry_1\ : std_logic;
signal \alogicunit.un1_a_1_cry_2_THRU_CO\ : std_logic;
signal \alogicunit.un1_a_1_cry_2\ : std_logic;
signal \alogicunit.un1_a_1_cry_3\ : std_logic;
signal \alogicunit.result_RNO_0Z0Z_5\ : std_logic;
signal \alogicunit.un1_a_1_cry_4\ : std_logic;
signal \alogicunit.un1_a_1_cry_5\ : std_logic;
signal \alogicunit.N_95_1\ : std_logic;
signal \alogicunit.un1_a_1_cry_6\ : std_logic;
signal left_3 : std_logic;
signal \alogicunit.m26_l_fxZ0Z_0\ : std_logic;
signal \un1_click13_1_sn_cascade_\ : std_logic;
signal \sevsegr_RNO_0Z0Z_2\ : std_logic;
signal \sevsegr_RNO_0Z0Z_1\ : std_logic;
signal \r_SwitchZ0Z_3\ : std_logic;
signal \alogicunit.m26_l_fxZ0\ : std_logic;
signal \sevsegl_RNO_0Z0Z_1\ : std_logic;
signal \r_CountZ0Z_3\ : std_logic;
signal \sevsegl_RNO_0Z0Z_3\ : std_logic;
signal \alogicunit.result24\ : std_logic;
signal \alogicunit.result24_cascade_\ : std_logic;
signal \alogicunit.un1_a_1_axb_3\ : std_logic;
signal \alogicunit.N_51\ : std_logic;
signal cu1_track_ns_3 : std_logic;
signal \N_28\ : std_logic;
signal \alogicunit.N_41\ : std_logic;
signal \alogicunit.N_41_cascade_\ : std_logic;
signal \track_RNI9MAL_0_1\ : std_logic;
signal \r_CountZ0Z_1\ : std_logic;
signal \r_CountZ0Z_0\ : std_logic;
signal \r_CountZ0Z_2\ : std_logic;
signal \Instance2.r_Count13_8_0_cascade_\ : std_logic;
signal \Instance2.un1_r_Count_10lt11_0_cascade_\ : std_logic;
signal \Instance2.r_Count13_12\ : std_logic;
signal \Instance2.r_Count13_13_cascade_\ : std_logic;
signal \Instance2.un1_r_Count_10lto11_1\ : std_logic;
signal \Instance2.r_Count13_10\ : std_logic;
signal \Instance2.r_Count13_7\ : std_logic;
signal \alogicunit.N_90\ : std_logic;
signal \Instance2.r_Count13_4\ : std_logic;
signal click13 : std_logic;
signal \alogicunit.N_49\ : std_logic;
signal \r_SwitchZ0Z_2\ : std_logic;
signal \r_SwitchZ0Z_4\ : std_logic;
signal \Instance2.click14_sn_cascade_\ : std_logic;
signal un1_click13_1_sn : std_logic;
signal \Instance2_un1_click13_3_1\ : std_logic;
signal \alogicunit.result_RNO_0Z0Z_4\ : std_logic;
signal left_0 : std_logic;
signal \alogicunit.N_50\ : std_logic;
signal \alogicunit.result_RNO_0Z0Z_6\ : std_logic;
signal left_2 : std_logic;
signal \alogicunit.un1_a_1_cry_1_c_invZ0\ : std_logic;
signal \alogicunit.N_102\ : std_logic;
signal \r_HexEncode_i_0_4\ : std_logic;
signal \alogicunit.N_35\ : std_logic;
signal \alogicunit.result24_iZ0\ : std_logic;
signal current_state_0 : std_logic;
signal current_state_1 : std_logic;
signal current_state_2 : std_logic;
signal current_state_3 : std_logic;
signal \clickZ0Z1\ : std_logic;
signal \Instance2.un1_r_Count_10lto17_1\ : std_logic;
signal \w_Switch_2\ : std_logic;
signal \i_Switch_2_c\ : std_logic;
signal \Instance2.un1_r_Count_10lt17\ : std_logic;
signal \Instance2.r_Count12_i\ : std_logic;
signal \bfn_6_7_0_\ : std_logic;
signal \Instance4.r_Count_2_cry_1\ : std_logic;
signal \Instance4.r_Count_2_cry_2\ : std_logic;
signal \Instance4.r_Count_2_cry_3\ : std_logic;
signal \Instance4.r_Count_2_cry_4\ : std_logic;
signal \Instance4.r_Count_2_cry_5\ : std_logic;
signal \Instance4.r_Count_2_cry_6\ : std_logic;
signal \Instance4.r_Count_2_cry_7\ : std_logic;
signal \Instance4.r_Count_2_cry_8\ : std_logic;
signal \bfn_6_8_0_\ : std_logic;
signal \Instance4.r_Count_2_cry_9\ : std_logic;
signal \Instance4.r_Count_2_cry_10\ : std_logic;
signal \Instance4.r_Count_2_cry_11\ : std_logic;
signal \Instance4.r_Count_2_cry_12\ : std_logic;
signal \Instance4.r_Count_2_cry_13\ : std_logic;
signal \Instance4.r_Count_2_cry_14\ : std_logic;
signal \Instance4.r_Count_2_cry_15\ : std_logic;
signal \Instance4.r_Count_2_cry_16\ : std_logic;
signal \bfn_6_9_0_\ : std_logic;
signal \Instance4.r_Count12_i_g\ : std_logic;
signal \bfn_6_10_0_\ : std_logic;
signal \Instance2.r_Count_0_2\ : std_logic;
signal \Instance2.r_Count_2_cry_1\ : std_logic;
signal \Instance2.r_Count_0_3\ : std_logic;
signal \Instance2.r_Count_2_cry_2\ : std_logic;
signal \Instance2.r_CountZ0Z_4\ : std_logic;
signal \Instance2.r_Count_2_cry_3\ : std_logic;
signal \Instance2.r_CountZ0Z_5\ : std_logic;
signal \Instance2.r_Count_2_cry_4\ : std_logic;
signal \Instance2.r_CountZ0Z_6\ : std_logic;
signal \Instance2.r_Count_2_cry_5\ : std_logic;
signal \Instance2.r_CountZ0Z_7\ : std_logic;
signal \Instance2.r_Count_2_cry_6\ : std_logic;
signal \Instance2.r_CountZ0Z_8\ : std_logic;
signal \Instance2.r_Count_2_cry_7\ : std_logic;
signal \Instance2.r_Count_2_cry_8\ : std_logic;
signal \Instance2.r_CountZ0Z_9\ : std_logic;
signal \bfn_6_11_0_\ : std_logic;
signal \Instance2.r_CountZ0Z_10\ : std_logic;
signal \Instance2.r_Count_2_cry_9\ : std_logic;
signal \Instance2.r_CountZ0Z_11\ : std_logic;
signal \Instance2.r_Count_2_cry_10\ : std_logic;
signal \Instance2.r_CountZ0Z_12\ : std_logic;
signal \Instance2.r_Count_2_cry_11\ : std_logic;
signal \Instance2.r_CountZ0Z_13\ : std_logic;
signal \Instance2.r_Count_2_cry_12\ : std_logic;
signal \Instance2.r_CountZ0Z_14\ : std_logic;
signal \Instance2.r_Count_2_cry_13\ : std_logic;
signal \Instance2.r_CountZ0Z_15\ : std_logic;
signal \Instance2.r_Count_2_cry_14\ : std_logic;
signal \Instance2.r_CountZ0Z_16\ : std_logic;
signal \Instance2.r_Count_2_cry_15\ : std_logic;
signal \Instance2.r_Count_2_cry_16\ : std_logic;
signal \bfn_6_12_0_\ : std_logic;
signal \Instance2.r_CountZ0Z_17\ : std_logic;
signal \Instance2.r_Count_0_0\ : std_logic;
signal \Instance2.r_Count_0_1\ : std_logic;
signal \Instance2.r_Count12_i_g\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \r_HexEncode_i_0_3\ : std_logic;
signal \sevseglZ0Z_2\ : std_logic;
signal \sevseglZ0Z_1\ : std_logic;
signal \sevseglZ0Z_3\ : std_logic;
signal \sevseglZ0Z_0\ : std_logic;
signal \r_HexEncode_i_0_2\ : std_logic;
signal \Instance4.r_CountZ0Z_1\ : std_logic;
signal \Instance4.r_CountZ0Z_2\ : std_logic;
signal \Instance4.r_CountZ0Z_3\ : std_logic;
signal \Instance4.r_CountZ0Z_4\ : std_logic;
signal \Instance4.r_CountZ0Z_7\ : std_logic;
signal \Instance4.r_CountZ0Z_0\ : std_logic;
signal \Instance4.r_Count13_8_0_cascade_\ : std_logic;
signal \Instance4.r_CountZ0Z_5\ : std_logic;
signal \Instance4.r_Count13_7\ : std_logic;
signal \Instance4.r_Count13_13_cascade_\ : std_logic;
signal \Instance4.r_Count13_12\ : std_logic;
signal \Instance4.r_CountZ0Z_14\ : std_logic;
signal \Instance4.r_CountZ0Z_17\ : std_logic;
signal \Instance4.r_Count13_4\ : std_logic;
signal \Instance4.r_CountZ0Z_11\ : std_logic;
signal \Instance4.r_CountZ0Z_10\ : std_logic;
signal \Instance4.r_CountZ0Z_9\ : std_logic;
signal \Instance4.r_CountZ0Z_13\ : std_logic;
signal \Instance4.r_CountZ0Z_12\ : std_logic;
signal \Instance4.un1_r_Count_10lto11_1_cascade_\ : std_logic;
signal \Instance4.un1_r_Count_10lt11_0\ : std_logic;
signal \i_Switch_4_c\ : std_logic;
signal \w_Switch_4\ : std_logic;
signal \Instance4.un1_r_Count_10lt17_cascade_\ : std_logic;
signal \Instance4.un1_r_Count_10lto17_1\ : std_logic;
signal \Instance4.r_Count12_i\ : std_logic;
signal \Instance4.r_CountZ0Z_8\ : std_logic;
signal \Instance4.r_CountZ0Z_15\ : std_logic;
signal \Instance4.r_CountZ0Z_16\ : std_logic;
signal \Instance4.r_CountZ0Z_6\ : std_logic;
signal \Instance4.r_Count13_10\ : std_logic;
signal \w_Switch_3\ : std_logic;
signal \i_Switch_3_c\ : std_logic;
signal \Instance3.un1_r_Count_10lt17_cascade_\ : std_logic;
signal \Instance3.r_Count12_i\ : std_logic;
signal \Instance3.r_Count13_8_0_cascade_\ : std_logic;
signal \Instance3.r_Count13_12\ : std_logic;
signal \Instance3.un1_r_Count_10lt11_0\ : std_logic;
signal \Instance3.un1_r_Count_10lto11_1\ : std_logic;
signal \Instance3.r_Count13_4\ : std_logic;
signal \Instance3.r_Count13_7_cascade_\ : std_logic;
signal \Instance3.r_Count13_13\ : std_logic;
signal \Instance3.r_Count13_10\ : std_logic;
signal \Instance3.un1_r_Count_10lto17_1\ : std_logic;
signal negative : std_logic;
signal \o_LED_1_c\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \Instance3.r_CountZ0Z_2\ : std_logic;
signal \Instance3.r_Count_2_cry_1\ : std_logic;
signal \Instance3.r_CountZ0Z_3\ : std_logic;
signal \Instance3.r_Count_2_cry_2\ : std_logic;
signal \Instance3.r_CountZ0Z_4\ : std_logic;
signal \Instance3.r_Count_2_cry_3\ : std_logic;
signal \Instance3.r_CountZ0Z_5\ : std_logic;
signal \Instance3.r_Count_2_cry_4\ : std_logic;
signal \Instance3.r_CountZ0Z_6\ : std_logic;
signal \Instance3.r_Count_2_cry_5\ : std_logic;
signal \Instance3.r_CountZ0Z_7\ : std_logic;
signal \Instance3.r_Count_2_cry_6\ : std_logic;
signal \Instance3.r_CountZ0Z_8\ : std_logic;
signal \Instance3.r_Count_2_cry_7\ : std_logic;
signal \Instance3.r_Count_2_cry_8\ : std_logic;
signal \Instance3.r_CountZ0Z_9\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal \Instance3.r_CountZ0Z_10\ : std_logic;
signal \Instance3.r_Count_2_cry_9\ : std_logic;
signal \Instance3.r_CountZ0Z_11\ : std_logic;
signal \Instance3.r_Count_2_cry_10\ : std_logic;
signal \Instance3.r_CountZ0Z_12\ : std_logic;
signal \Instance3.r_Count_2_cry_11\ : std_logic;
signal \Instance3.r_CountZ0Z_13\ : std_logic;
signal \Instance3.r_Count_2_cry_12\ : std_logic;
signal \Instance3.r_CountZ0Z_14\ : std_logic;
signal \Instance3.r_Count_2_cry_13\ : std_logic;
signal \Instance3.r_CountZ0Z_15\ : std_logic;
signal \Instance3.r_Count_2_cry_14\ : std_logic;
signal \Instance3.r_CountZ0Z_16\ : std_logic;
signal \Instance3.r_Count_2_cry_15\ : std_logic;
signal \Instance3.r_Count_2_cry_16\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \Instance3.r_CountZ0Z_17\ : std_logic;
signal \Instance3.r_CountZ0Z_0\ : std_logic;
signal \Instance3.r_CountZ0Z_1\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \i_Clk_c_g\ : std_logic;
signal \Instance3.r_Count12_i_g\ : std_logic;

signal \i_Clk_wire\ : std_logic;
signal \o_Segment2_F_wire\ : std_logic;
signal \o_LED_1_wire\ : std_logic;
signal \o_Segment1_G_wire\ : std_logic;
signal \i_Switch_4_wire\ : std_logic;
signal \i_Switch_1_wire\ : std_logic;
signal \o_Segment1_B_wire\ : std_logic;
signal \i_Switch_3_wire\ : std_logic;
signal \o_Segment1_E_wire\ : std_logic;
signal \o_LED_2_wire\ : std_logic;
signal \o_Segment2_E_wire\ : std_logic;
signal \o_Segment2_C_wire\ : std_logic;
signal \o_LED_4_wire\ : std_logic;
signal \o_Segment1_A_wire\ : std_logic;
signal \i_Switch_2_wire\ : std_logic;
signal \o_Segment2_B_wire\ : std_logic;
signal \o_Segment1_C_wire\ : std_logic;
signal \o_Segment1_D_wire\ : std_logic;
signal \o_Segment1_F_wire\ : std_logic;
signal \o_LED_3_wire\ : std_logic;
signal \o_Segment2_A_wire\ : std_logic;
signal \o_Segment2_G_wire\ : std_logic;
signal \o_Segment2_D_wire\ : std_logic;

begin
    \i_Clk_wire\ <= i_Clk;
    o_Segment2_F <= \o_Segment2_F_wire\;
    o_LED_1 <= \o_LED_1_wire\;
    o_Segment1_G <= \o_Segment1_G_wire\;
    \i_Switch_4_wire\ <= i_Switch_4;
    \i_Switch_1_wire\ <= i_Switch_1;
    o_Segment1_B <= \o_Segment1_B_wire\;
    \i_Switch_3_wire\ <= i_Switch_3;
    o_Segment1_E <= \o_Segment1_E_wire\;
    o_LED_2 <= \o_LED_2_wire\;
    o_Segment2_E <= \o_Segment2_E_wire\;
    o_Segment2_C <= \o_Segment2_C_wire\;
    o_LED_4 <= \o_LED_4_wire\;
    o_Segment1_A <= \o_Segment1_A_wire\;
    \i_Switch_2_wire\ <= i_Switch_2;
    o_Segment2_B <= \o_Segment2_B_wire\;
    o_Segment1_C <= \o_Segment1_C_wire\;
    o_Segment1_D <= \o_Segment1_D_wire\;
    o_Segment1_F <= \o_Segment1_F_wire\;
    o_LED_3 <= \o_LED_3_wire\;
    o_Segment2_A <= \o_Segment2_A_wire\;
    o_Segment2_G <= \o_Segment2_G_wire\;
    o_Segment2_D <= \o_Segment2_D_wire\;

    \i_Clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__7468\,
            GLOBALBUFFEROUTPUT => \i_Clk_c_g\
        );

    \i_Clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7470\,
            DIN => \N__7469\,
            DOUT => \N__7468\,
            PACKAGEPIN => \i_Clk_wire\
        );

    \i_Clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7470\,
            PADOUT => \N__7469\,
            PADIN => \N__7468\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_Segment2_F_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7459\,
            DIN => \N__7458\,
            DOUT => \N__7457\,
            PACKAGEPIN => \o_Segment2_F_wire\
        );

    \o_Segment2_F_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7459\,
            PADOUT => \N__7458\,
            PADIN => \N__7457\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3111\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_LED_1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7450\,
            DIN => \N__7449\,
            DOUT => \N__7448\,
            PACKAGEPIN => \o_LED_1_wire\
        );

    \o_LED_1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7450\,
            PADOUT => \N__7449\,
            PADIN => \N__7448\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6759\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_Segment1_G_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7441\,
            DIN => \N__7440\,
            DOUT => \N__7439\,
            PACKAGEPIN => \o_Segment1_G_wire\
        );

    \o_Segment1_G_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7441\,
            PADOUT => \N__7440\,
            PADIN => \N__7439\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3240\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \i_Switch_4_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7432\,
            DIN => \N__7431\,
            DOUT => \N__7430\,
            PACKAGEPIN => \i_Switch_4_wire\
        );

    \i_Switch_4_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7432\,
            PADOUT => \N__7431\,
            PADIN => \N__7430\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \i_Switch_4_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \i_Switch_1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7423\,
            DIN => \N__7422\,
            DOUT => \N__7421\,
            PACKAGEPIN => \i_Switch_1_wire\
        );

    \i_Switch_1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7423\,
            PADOUT => \N__7422\,
            PADIN => \N__7421\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \i_Switch_1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_Segment1_B_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7414\,
            DIN => \N__7413\,
            DOUT => \N__7412\,
            PACKAGEPIN => \o_Segment1_B_wire\
        );

    \o_Segment1_B_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7414\,
            PADOUT => \N__7413\,
            PADIN => \N__7412\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3105\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \i_Switch_3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7405\,
            DIN => \N__7404\,
            DOUT => \N__7403\,
            PACKAGEPIN => \i_Switch_3_wire\
        );

    \i_Switch_3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7405\,
            PADOUT => \N__7404\,
            PADIN => \N__7403\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \i_Switch_3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_Segment1_E_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7396\,
            DIN => \N__7395\,
            DOUT => \N__7394\,
            PACKAGEPIN => \o_Segment1_E_wire\
        );

    \o_Segment1_E_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7396\,
            PADOUT => \N__7395\,
            PADIN => \N__7394\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5892\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_LED_2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7387\,
            DIN => \N__7386\,
            DOUT => \N__7385\,
            PACKAGEPIN => \o_LED_2_wire\
        );

    \o_LED_2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7387\,
            PADOUT => \N__7386\,
            PADIN => \N__7385\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6757\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_Segment2_E_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7378\,
            DIN => \N__7377\,
            DOUT => \N__7376\,
            PACKAGEPIN => \o_Segment2_E_wire\
        );

    \o_Segment2_E_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7378\,
            PADOUT => \N__7377\,
            PADIN => \N__7376\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3804\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_Segment2_C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7369\,
            DIN => \N__7368\,
            DOUT => \N__7367\,
            PACKAGEPIN => \o_Segment2_C_wire\
        );

    \o_Segment2_C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7369\,
            PADOUT => \N__7368\,
            PADIN => \N__7367\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3825\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_LED_4_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7360\,
            DIN => \N__7359\,
            DOUT => \N__7358\,
            PACKAGEPIN => \o_LED_4_wire\
        );

    \o_LED_4_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7360\,
            PADOUT => \N__7359\,
            PADIN => \N__7358\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6747\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_Segment1_A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7351\,
            DIN => \N__7350\,
            DOUT => \N__7349\,
            PACKAGEPIN => \o_Segment1_A_wire\
        );

    \o_Segment1_A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7351\,
            PADOUT => \N__7350\,
            PADIN => \N__7349\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3117\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \i_Switch_2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7342\,
            DIN => \N__7341\,
            DOUT => \N__7340\,
            PACKAGEPIN => \i_Switch_2_wire\
        );

    \i_Switch_2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7342\,
            PADOUT => \N__7341\,
            PADIN => \N__7340\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \i_Switch_2_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_Segment2_B_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7333\,
            DIN => \N__7332\,
            DOUT => \N__7331\,
            PACKAGEPIN => \o_Segment2_B_wire\
        );

    \o_Segment2_B_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7333\,
            PADOUT => \N__7332\,
            PADIN => \N__7331\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3621\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_Segment1_C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7324\,
            DIN => \N__7323\,
            DOUT => \N__7322\,
            PACKAGEPIN => \o_Segment1_C_wire\
        );

    \o_Segment1_C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7324\,
            PADOUT => \N__7323\,
            PADIN => \N__7322\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5415\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_Segment1_D_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7315\,
            DIN => \N__7314\,
            DOUT => \N__7313\,
            PACKAGEPIN => \o_Segment1_D_wire\
        );

    \o_Segment1_D_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7315\,
            PADOUT => \N__7314\,
            PADIN => \N__7313\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6087\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_Segment1_F_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7306\,
            DIN => \N__7305\,
            DOUT => \N__7304\,
            PACKAGEPIN => \o_Segment1_F_wire\
        );

    \o_Segment1_F_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7306\,
            PADOUT => \N__7305\,
            PADIN => \N__7304\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3234\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_LED_3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7297\,
            DIN => \N__7296\,
            DOUT => \N__7295\,
            PACKAGEPIN => \o_LED_3_wire\
        );

    \o_LED_3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7297\,
            PADOUT => \N__7296\,
            PADIN => \N__7295\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6758\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_Segment2_A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7288\,
            DIN => \N__7287\,
            DOUT => \N__7286\,
            PACKAGEPIN => \o_Segment2_A_wire\
        );

    \o_Segment2_A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7288\,
            PADOUT => \N__7287\,
            PADIN => \N__7286\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3228\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_Segment2_G_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7279\,
            DIN => \N__7278\,
            DOUT => \N__7277\,
            PACKAGEPIN => \o_Segment2_G_wire\
        );

    \o_Segment2_G_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7279\,
            PADOUT => \N__7278\,
            PADIN => \N__7277\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3819\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_Segment2_D_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7270\,
            DIN => \N__7269\,
            DOUT => \N__7268\,
            PACKAGEPIN => \o_Segment2_D_wire\
        );

    \o_Segment2_D_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7270\,
            PADOUT => \N__7269\,
            PADIN => \N__7268\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3792\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1682\ : CascadeMux
    port map (
            O => \N__7251\,
            I => \N__7246\
        );

    \I__1681\ : InMux
    port map (
            O => \N__7250\,
            I => \N__7243\
        );

    \I__1680\ : InMux
    port map (
            O => \N__7249\,
            I => \N__7238\
        );

    \I__1679\ : InMux
    port map (
            O => \N__7246\,
            I => \N__7238\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__7243\,
            I => \Instance3.r_CountZ0Z_14\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__7238\,
            I => \Instance3.r_CountZ0Z_14\
        );

    \I__1676\ : InMux
    port map (
            O => \N__7233\,
            I => \Instance3.r_Count_2_cry_13\
        );

    \I__1675\ : CascadeMux
    port map (
            O => \N__7230\,
            I => \N__7226\
        );

    \I__1674\ : InMux
    port map (
            O => \N__7229\,
            I => \N__7222\
        );

    \I__1673\ : InMux
    port map (
            O => \N__7226\,
            I => \N__7219\
        );

    \I__1672\ : InMux
    port map (
            O => \N__7225\,
            I => \N__7216\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__7222\,
            I => \Instance3.r_CountZ0Z_15\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__7219\,
            I => \Instance3.r_CountZ0Z_15\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__7216\,
            I => \Instance3.r_CountZ0Z_15\
        );

    \I__1668\ : InMux
    port map (
            O => \N__7209\,
            I => \Instance3.r_Count_2_cry_14\
        );

    \I__1667\ : InMux
    port map (
            O => \N__7206\,
            I => \N__7201\
        );

    \I__1666\ : InMux
    port map (
            O => \N__7205\,
            I => \N__7198\
        );

    \I__1665\ : InMux
    port map (
            O => \N__7204\,
            I => \N__7195\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__7201\,
            I => \Instance3.r_CountZ0Z_16\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__7198\,
            I => \Instance3.r_CountZ0Z_16\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__7195\,
            I => \Instance3.r_CountZ0Z_16\
        );

    \I__1661\ : InMux
    port map (
            O => \N__7188\,
            I => \Instance3.r_Count_2_cry_15\
        );

    \I__1660\ : InMux
    port map (
            O => \N__7185\,
            I => \bfn_8_11_0_\
        );

    \I__1659\ : InMux
    port map (
            O => \N__7182\,
            I => \N__7177\
        );

    \I__1658\ : InMux
    port map (
            O => \N__7181\,
            I => \N__7172\
        );

    \I__1657\ : InMux
    port map (
            O => \N__7180\,
            I => \N__7172\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__7177\,
            I => \Instance3.r_CountZ0Z_17\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__7172\,
            I => \Instance3.r_CountZ0Z_17\
        );

    \I__1654\ : InMux
    port map (
            O => \N__7167\,
            I => \N__7164\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__7164\,
            I => \N__7158\
        );

    \I__1652\ : CascadeMux
    port map (
            O => \N__7163\,
            I => \N__7155\
        );

    \I__1651\ : InMux
    port map (
            O => \N__7162\,
            I => \N__7150\
        );

    \I__1650\ : InMux
    port map (
            O => \N__7161\,
            I => \N__7150\
        );

    \I__1649\ : Span4Mux_v
    port map (
            O => \N__7158\,
            I => \N__7147\
        );

    \I__1648\ : InMux
    port map (
            O => \N__7155\,
            I => \N__7144\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__7150\,
            I => \Instance3.r_CountZ0Z_0\
        );

    \I__1646\ : Odrv4
    port map (
            O => \N__7147\,
            I => \Instance3.r_CountZ0Z_0\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__7144\,
            I => \Instance3.r_CountZ0Z_0\
        );

    \I__1644\ : InMux
    port map (
            O => \N__7137\,
            I => \N__7132\
        );

    \I__1643\ : InMux
    port map (
            O => \N__7136\,
            I => \N__7129\
        );

    \I__1642\ : InMux
    port map (
            O => \N__7135\,
            I => \N__7126\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__7132\,
            I => \N__7123\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__7129\,
            I => \Instance3.r_CountZ0Z_1\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__7126\,
            I => \Instance3.r_CountZ0Z_1\
        );

    \I__1638\ : Odrv4
    port map (
            O => \N__7123\,
            I => \Instance3.r_CountZ0Z_1\
        );

    \I__1637\ : ClkMux
    port map (
            O => \N__7116\,
            I => \N__7008\
        );

    \I__1636\ : ClkMux
    port map (
            O => \N__7115\,
            I => \N__7008\
        );

    \I__1635\ : ClkMux
    port map (
            O => \N__7114\,
            I => \N__7008\
        );

    \I__1634\ : ClkMux
    port map (
            O => \N__7113\,
            I => \N__7008\
        );

    \I__1633\ : ClkMux
    port map (
            O => \N__7112\,
            I => \N__7008\
        );

    \I__1632\ : ClkMux
    port map (
            O => \N__7111\,
            I => \N__7008\
        );

    \I__1631\ : ClkMux
    port map (
            O => \N__7110\,
            I => \N__7008\
        );

    \I__1630\ : ClkMux
    port map (
            O => \N__7109\,
            I => \N__7008\
        );

    \I__1629\ : ClkMux
    port map (
            O => \N__7108\,
            I => \N__7008\
        );

    \I__1628\ : ClkMux
    port map (
            O => \N__7107\,
            I => \N__7008\
        );

    \I__1627\ : ClkMux
    port map (
            O => \N__7106\,
            I => \N__7008\
        );

    \I__1626\ : ClkMux
    port map (
            O => \N__7105\,
            I => \N__7008\
        );

    \I__1625\ : ClkMux
    port map (
            O => \N__7104\,
            I => \N__7008\
        );

    \I__1624\ : ClkMux
    port map (
            O => \N__7103\,
            I => \N__7008\
        );

    \I__1623\ : ClkMux
    port map (
            O => \N__7102\,
            I => \N__7008\
        );

    \I__1622\ : ClkMux
    port map (
            O => \N__7101\,
            I => \N__7008\
        );

    \I__1621\ : ClkMux
    port map (
            O => \N__7100\,
            I => \N__7008\
        );

    \I__1620\ : ClkMux
    port map (
            O => \N__7099\,
            I => \N__7008\
        );

    \I__1619\ : ClkMux
    port map (
            O => \N__7098\,
            I => \N__7008\
        );

    \I__1618\ : ClkMux
    port map (
            O => \N__7097\,
            I => \N__7008\
        );

    \I__1617\ : ClkMux
    port map (
            O => \N__7096\,
            I => \N__7008\
        );

    \I__1616\ : ClkMux
    port map (
            O => \N__7095\,
            I => \N__7008\
        );

    \I__1615\ : ClkMux
    port map (
            O => \N__7094\,
            I => \N__7008\
        );

    \I__1614\ : ClkMux
    port map (
            O => \N__7093\,
            I => \N__7008\
        );

    \I__1613\ : ClkMux
    port map (
            O => \N__7092\,
            I => \N__7008\
        );

    \I__1612\ : ClkMux
    port map (
            O => \N__7091\,
            I => \N__7008\
        );

    \I__1611\ : ClkMux
    port map (
            O => \N__7090\,
            I => \N__7008\
        );

    \I__1610\ : ClkMux
    port map (
            O => \N__7089\,
            I => \N__7008\
        );

    \I__1609\ : ClkMux
    port map (
            O => \N__7088\,
            I => \N__7008\
        );

    \I__1608\ : ClkMux
    port map (
            O => \N__7087\,
            I => \N__7008\
        );

    \I__1607\ : ClkMux
    port map (
            O => \N__7086\,
            I => \N__7008\
        );

    \I__1606\ : ClkMux
    port map (
            O => \N__7085\,
            I => \N__7008\
        );

    \I__1605\ : ClkMux
    port map (
            O => \N__7084\,
            I => \N__7008\
        );

    \I__1604\ : ClkMux
    port map (
            O => \N__7083\,
            I => \N__7008\
        );

    \I__1603\ : ClkMux
    port map (
            O => \N__7082\,
            I => \N__7008\
        );

    \I__1602\ : ClkMux
    port map (
            O => \N__7081\,
            I => \N__7008\
        );

    \I__1601\ : GlobalMux
    port map (
            O => \N__7008\,
            I => \N__7005\
        );

    \I__1600\ : gio2CtrlBuf
    port map (
            O => \N__7005\,
            I => \i_Clk_c_g\
        );

    \I__1599\ : SRMux
    port map (
            O => \N__7002\,
            I => \N__6990\
        );

    \I__1598\ : SRMux
    port map (
            O => \N__7001\,
            I => \N__6990\
        );

    \I__1597\ : SRMux
    port map (
            O => \N__7000\,
            I => \N__6990\
        );

    \I__1596\ : SRMux
    port map (
            O => \N__6999\,
            I => \N__6990\
        );

    \I__1595\ : GlobalMux
    port map (
            O => \N__6990\,
            I => \N__6987\
        );

    \I__1594\ : gio2CtrlBuf
    port map (
            O => \N__6987\,
            I => \Instance3.r_Count12_i_g\
        );

    \I__1593\ : InMux
    port map (
            O => \N__6984\,
            I => \Instance3.r_Count_2_cry_4\
        );

    \I__1592\ : CascadeMux
    port map (
            O => \N__6981\,
            I => \N__6976\
        );

    \I__1591\ : InMux
    port map (
            O => \N__6980\,
            I => \N__6973\
        );

    \I__1590\ : InMux
    port map (
            O => \N__6979\,
            I => \N__6970\
        );

    \I__1589\ : InMux
    port map (
            O => \N__6976\,
            I => \N__6967\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__6973\,
            I => \Instance3.r_CountZ0Z_6\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__6970\,
            I => \Instance3.r_CountZ0Z_6\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__6967\,
            I => \Instance3.r_CountZ0Z_6\
        );

    \I__1585\ : InMux
    port map (
            O => \N__6960\,
            I => \Instance3.r_Count_2_cry_5\
        );

    \I__1584\ : InMux
    port map (
            O => \N__6957\,
            I => \N__6952\
        );

    \I__1583\ : InMux
    port map (
            O => \N__6956\,
            I => \N__6947\
        );

    \I__1582\ : InMux
    port map (
            O => \N__6955\,
            I => \N__6947\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__6952\,
            I => \Instance3.r_CountZ0Z_7\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__6947\,
            I => \Instance3.r_CountZ0Z_7\
        );

    \I__1579\ : InMux
    port map (
            O => \N__6942\,
            I => \Instance3.r_Count_2_cry_6\
        );

    \I__1578\ : InMux
    port map (
            O => \N__6939\,
            I => \N__6934\
        );

    \I__1577\ : InMux
    port map (
            O => \N__6938\,
            I => \N__6931\
        );

    \I__1576\ : InMux
    port map (
            O => \N__6937\,
            I => \N__6928\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__6934\,
            I => \Instance3.r_CountZ0Z_8\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__6931\,
            I => \Instance3.r_CountZ0Z_8\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__6928\,
            I => \Instance3.r_CountZ0Z_8\
        );

    \I__1572\ : InMux
    port map (
            O => \N__6921\,
            I => \Instance3.r_Count_2_cry_7\
        );

    \I__1571\ : InMux
    port map (
            O => \N__6918\,
            I => \N__6913\
        );

    \I__1570\ : InMux
    port map (
            O => \N__6917\,
            I => \N__6910\
        );

    \I__1569\ : InMux
    port map (
            O => \N__6916\,
            I => \N__6907\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__6913\,
            I => \Instance3.r_CountZ0Z_9\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__6910\,
            I => \Instance3.r_CountZ0Z_9\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__6907\,
            I => \Instance3.r_CountZ0Z_9\
        );

    \I__1565\ : InMux
    port map (
            O => \N__6900\,
            I => \bfn_8_10_0_\
        );

    \I__1564\ : CascadeMux
    port map (
            O => \N__6897\,
            I => \N__6894\
        );

    \I__1563\ : InMux
    port map (
            O => \N__6894\,
            I => \N__6889\
        );

    \I__1562\ : InMux
    port map (
            O => \N__6893\,
            I => \N__6886\
        );

    \I__1561\ : InMux
    port map (
            O => \N__6892\,
            I => \N__6883\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__6889\,
            I => \N__6880\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__6886\,
            I => \Instance3.r_CountZ0Z_10\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__6883\,
            I => \Instance3.r_CountZ0Z_10\
        );

    \I__1557\ : Odrv4
    port map (
            O => \N__6880\,
            I => \Instance3.r_CountZ0Z_10\
        );

    \I__1556\ : InMux
    port map (
            O => \N__6873\,
            I => \Instance3.r_Count_2_cry_9\
        );

    \I__1555\ : InMux
    port map (
            O => \N__6870\,
            I => \N__6865\
        );

    \I__1554\ : InMux
    port map (
            O => \N__6869\,
            I => \N__6862\
        );

    \I__1553\ : InMux
    port map (
            O => \N__6868\,
            I => \N__6859\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__6865\,
            I => \N__6856\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__6862\,
            I => \Instance3.r_CountZ0Z_11\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__6859\,
            I => \Instance3.r_CountZ0Z_11\
        );

    \I__1549\ : Odrv4
    port map (
            O => \N__6856\,
            I => \Instance3.r_CountZ0Z_11\
        );

    \I__1548\ : InMux
    port map (
            O => \N__6849\,
            I => \Instance3.r_Count_2_cry_10\
        );

    \I__1547\ : CascadeMux
    port map (
            O => \N__6846\,
            I => \N__6843\
        );

    \I__1546\ : InMux
    port map (
            O => \N__6843\,
            I => \N__6838\
        );

    \I__1545\ : InMux
    port map (
            O => \N__6842\,
            I => \N__6835\
        );

    \I__1544\ : InMux
    port map (
            O => \N__6841\,
            I => \N__6832\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__6838\,
            I => \N__6829\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__6835\,
            I => \Instance3.r_CountZ0Z_12\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__6832\,
            I => \Instance3.r_CountZ0Z_12\
        );

    \I__1540\ : Odrv4
    port map (
            O => \N__6829\,
            I => \Instance3.r_CountZ0Z_12\
        );

    \I__1539\ : InMux
    port map (
            O => \N__6822\,
            I => \Instance3.r_Count_2_cry_11\
        );

    \I__1538\ : CascadeMux
    port map (
            O => \N__6819\,
            I => \N__6815\
        );

    \I__1537\ : InMux
    port map (
            O => \N__6818\,
            I => \N__6811\
        );

    \I__1536\ : InMux
    port map (
            O => \N__6815\,
            I => \N__6806\
        );

    \I__1535\ : InMux
    port map (
            O => \N__6814\,
            I => \N__6806\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__6811\,
            I => \Instance3.r_CountZ0Z_13\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__6806\,
            I => \Instance3.r_CountZ0Z_13\
        );

    \I__1532\ : InMux
    port map (
            O => \N__6801\,
            I => \Instance3.r_Count_2_cry_12\
        );

    \I__1531\ : CascadeMux
    port map (
            O => \N__6798\,
            I => \Instance3.r_Count13_7_cascade_\
        );

    \I__1530\ : InMux
    port map (
            O => \N__6795\,
            I => \N__6792\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__6792\,
            I => \N__6789\
        );

    \I__1528\ : Span4Mux_v
    port map (
            O => \N__6789\,
            I => \N__6786\
        );

    \I__1527\ : Odrv4
    port map (
            O => \N__6786\,
            I => \Instance3.r_Count13_13\
        );

    \I__1526\ : InMux
    port map (
            O => \N__6783\,
            I => \N__6780\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__6780\,
            I => \Instance3.r_Count13_10\
        );

    \I__1524\ : InMux
    port map (
            O => \N__6777\,
            I => \N__6774\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__6774\,
            I => \Instance3.un1_r_Count_10lto17_1\
        );

    \I__1522\ : InMux
    port map (
            O => \N__6771\,
            I => \N__6768\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__6768\,
            I => \N__6765\
        );

    \I__1520\ : Span4Mux_h
    port map (
            O => \N__6765\,
            I => \N__6762\
        );

    \I__1519\ : Odrv4
    port map (
            O => \N__6762\,
            I => negative
        );

    \I__1518\ : IoInMux
    port map (
            O => \N__6759\,
            I => \N__6754\
        );

    \I__1517\ : IoInMux
    port map (
            O => \N__6758\,
            I => \N__6751\
        );

    \I__1516\ : IoInMux
    port map (
            O => \N__6757\,
            I => \N__6748\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__6754\,
            I => \N__6744\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__6751\,
            I => \N__6739\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__6748\,
            I => \N__6739\
        );

    \I__1512\ : IoInMux
    port map (
            O => \N__6747\,
            I => \N__6736\
        );

    \I__1511\ : Span4Mux_s3_h
    port map (
            O => \N__6744\,
            I => \N__6733\
        );

    \I__1510\ : Span4Mux_s3_h
    port map (
            O => \N__6739\,
            I => \N__6730\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__6736\,
            I => \N__6727\
        );

    \I__1508\ : Odrv4
    port map (
            O => \N__6733\,
            I => \o_LED_1_c\
        );

    \I__1507\ : Odrv4
    port map (
            O => \N__6730\,
            I => \o_LED_1_c\
        );

    \I__1506\ : Odrv12
    port map (
            O => \N__6727\,
            I => \o_LED_1_c\
        );

    \I__1505\ : InMux
    port map (
            O => \N__6720\,
            I => \N__6716\
        );

    \I__1504\ : InMux
    port map (
            O => \N__6719\,
            I => \N__6713\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__6716\,
            I => \Instance3.r_CountZ0Z_2\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__6713\,
            I => \Instance3.r_CountZ0Z_2\
        );

    \I__1501\ : InMux
    port map (
            O => \N__6708\,
            I => \Instance3.r_Count_2_cry_1\
        );

    \I__1500\ : CascadeMux
    port map (
            O => \N__6705\,
            I => \N__6701\
        );

    \I__1499\ : InMux
    port map (
            O => \N__6704\,
            I => \N__6698\
        );

    \I__1498\ : InMux
    port map (
            O => \N__6701\,
            I => \N__6695\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__6698\,
            I => \Instance3.r_CountZ0Z_3\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__6695\,
            I => \Instance3.r_CountZ0Z_3\
        );

    \I__1495\ : InMux
    port map (
            O => \N__6690\,
            I => \Instance3.r_Count_2_cry_2\
        );

    \I__1494\ : InMux
    port map (
            O => \N__6687\,
            I => \N__6682\
        );

    \I__1493\ : InMux
    port map (
            O => \N__6686\,
            I => \N__6677\
        );

    \I__1492\ : InMux
    port map (
            O => \N__6685\,
            I => \N__6677\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__6682\,
            I => \Instance3.r_CountZ0Z_4\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__6677\,
            I => \Instance3.r_CountZ0Z_4\
        );

    \I__1489\ : InMux
    port map (
            O => \N__6672\,
            I => \Instance3.r_Count_2_cry_3\
        );

    \I__1488\ : InMux
    port map (
            O => \N__6669\,
            I => \N__6664\
        );

    \I__1487\ : InMux
    port map (
            O => \N__6668\,
            I => \N__6661\
        );

    \I__1486\ : InMux
    port map (
            O => \N__6667\,
            I => \N__6658\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__6664\,
            I => \N__6655\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__6661\,
            I => \Instance3.r_CountZ0Z_5\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__6658\,
            I => \Instance3.r_CountZ0Z_5\
        );

    \I__1482\ : Odrv4
    port map (
            O => \N__6655\,
            I => \Instance3.r_CountZ0Z_5\
        );

    \I__1481\ : InMux
    port map (
            O => \N__6648\,
            I => \N__6643\
        );

    \I__1480\ : InMux
    port map (
            O => \N__6647\,
            I => \N__6640\
        );

    \I__1479\ : InMux
    port map (
            O => \N__6646\,
            I => \N__6637\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__6643\,
            I => \Instance4.r_CountZ0Z_8\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__6640\,
            I => \Instance4.r_CountZ0Z_8\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__6637\,
            I => \Instance4.r_CountZ0Z_8\
        );

    \I__1475\ : InMux
    port map (
            O => \N__6630\,
            I => \N__6625\
        );

    \I__1474\ : InMux
    port map (
            O => \N__6629\,
            I => \N__6622\
        );

    \I__1473\ : InMux
    port map (
            O => \N__6628\,
            I => \N__6619\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__6625\,
            I => \Instance4.r_CountZ0Z_15\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__6622\,
            I => \Instance4.r_CountZ0Z_15\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__6619\,
            I => \Instance4.r_CountZ0Z_15\
        );

    \I__1469\ : CascadeMux
    port map (
            O => \N__6612\,
            I => \N__6608\
        );

    \I__1468\ : InMux
    port map (
            O => \N__6611\,
            I => \N__6604\
        );

    \I__1467\ : InMux
    port map (
            O => \N__6608\,
            I => \N__6599\
        );

    \I__1466\ : InMux
    port map (
            O => \N__6607\,
            I => \N__6599\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__6604\,
            I => \Instance4.r_CountZ0Z_16\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__6599\,
            I => \Instance4.r_CountZ0Z_16\
        );

    \I__1463\ : InMux
    port map (
            O => \N__6594\,
            I => \N__6589\
        );

    \I__1462\ : InMux
    port map (
            O => \N__6593\,
            I => \N__6586\
        );

    \I__1461\ : InMux
    port map (
            O => \N__6592\,
            I => \N__6583\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__6589\,
            I => \Instance4.r_CountZ0Z_6\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__6586\,
            I => \Instance4.r_CountZ0Z_6\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__6583\,
            I => \Instance4.r_CountZ0Z_6\
        );

    \I__1457\ : CascadeMux
    port map (
            O => \N__6576\,
            I => \N__6573\
        );

    \I__1456\ : InMux
    port map (
            O => \N__6573\,
            I => \N__6570\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__6570\,
            I => \Instance4.r_Count13_10\
        );

    \I__1454\ : InMux
    port map (
            O => \N__6567\,
            I => \N__6564\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__6564\,
            I => \N__6561\
        );

    \I__1452\ : Span4Mux_v
    port map (
            O => \N__6561\,
            I => \N__6557\
        );

    \I__1451\ : InMux
    port map (
            O => \N__6560\,
            I => \N__6552\
        );

    \I__1450\ : Span4Mux_h
    port map (
            O => \N__6557\,
            I => \N__6549\
        );

    \I__1449\ : InMux
    port map (
            O => \N__6556\,
            I => \N__6544\
        );

    \I__1448\ : InMux
    port map (
            O => \N__6555\,
            I => \N__6544\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__6552\,
            I => \w_Switch_3\
        );

    \I__1446\ : Odrv4
    port map (
            O => \N__6549\,
            I => \w_Switch_3\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__6544\,
            I => \w_Switch_3\
        );

    \I__1444\ : CascadeMux
    port map (
            O => \N__6537\,
            I => \N__6534\
        );

    \I__1443\ : InMux
    port map (
            O => \N__6534\,
            I => \N__6531\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__6531\,
            I => \N__6527\
        );

    \I__1441\ : InMux
    port map (
            O => \N__6530\,
            I => \N__6524\
        );

    \I__1440\ : Span4Mux_v
    port map (
            O => \N__6527\,
            I => \N__6521\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__6524\,
            I => \N__6518\
        );

    \I__1438\ : Span4Mux_h
    port map (
            O => \N__6521\,
            I => \N__6515\
        );

    \I__1437\ : Span4Mux_v
    port map (
            O => \N__6518\,
            I => \N__6512\
        );

    \I__1436\ : IoSpan4Mux
    port map (
            O => \N__6515\,
            I => \N__6509\
        );

    \I__1435\ : Span4Mux_h
    port map (
            O => \N__6512\,
            I => \N__6506\
        );

    \I__1434\ : Odrv4
    port map (
            O => \N__6509\,
            I => \i_Switch_3_c\
        );

    \I__1433\ : Odrv4
    port map (
            O => \N__6506\,
            I => \i_Switch_3_c\
        );

    \I__1432\ : CascadeMux
    port map (
            O => \N__6501\,
            I => \Instance3.un1_r_Count_10lt17_cascade_\
        );

    \I__1431\ : IoInMux
    port map (
            O => \N__6498\,
            I => \N__6495\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__6495\,
            I => \N__6492\
        );

    \I__1429\ : Odrv12
    port map (
            O => \N__6492\,
            I => \Instance3.r_Count12_i\
        );

    \I__1428\ : CascadeMux
    port map (
            O => \N__6489\,
            I => \Instance3.r_Count13_8_0_cascade_\
        );

    \I__1427\ : InMux
    port map (
            O => \N__6486\,
            I => \N__6483\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__6483\,
            I => \N__6480\
        );

    \I__1425\ : Span4Mux_h
    port map (
            O => \N__6480\,
            I => \N__6477\
        );

    \I__1424\ : Odrv4
    port map (
            O => \N__6477\,
            I => \Instance3.r_Count13_12\
        );

    \I__1423\ : InMux
    port map (
            O => \N__6474\,
            I => \N__6471\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__6471\,
            I => \Instance3.un1_r_Count_10lt11_0\
        );

    \I__1421\ : InMux
    port map (
            O => \N__6468\,
            I => \N__6465\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__6465\,
            I => \Instance3.un1_r_Count_10lto11_1\
        );

    \I__1419\ : InMux
    port map (
            O => \N__6462\,
            I => \N__6459\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__6459\,
            I => \Instance3.r_Count13_4\
        );

    \I__1417\ : CascadeMux
    port map (
            O => \N__6456\,
            I => \N__6450\
        );

    \I__1416\ : InMux
    port map (
            O => \N__6455\,
            I => \N__6445\
        );

    \I__1415\ : InMux
    port map (
            O => \N__6454\,
            I => \N__6445\
        );

    \I__1414\ : InMux
    port map (
            O => \N__6453\,
            I => \N__6442\
        );

    \I__1413\ : InMux
    port map (
            O => \N__6450\,
            I => \N__6439\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__6445\,
            I => \Instance4.r_CountZ0Z_0\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__6442\,
            I => \Instance4.r_CountZ0Z_0\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__6439\,
            I => \Instance4.r_CountZ0Z_0\
        );

    \I__1409\ : CascadeMux
    port map (
            O => \N__6432\,
            I => \Instance4.r_Count13_8_0_cascade_\
        );

    \I__1408\ : CascadeMux
    port map (
            O => \N__6429\,
            I => \N__6424\
        );

    \I__1407\ : InMux
    port map (
            O => \N__6428\,
            I => \N__6421\
        );

    \I__1406\ : InMux
    port map (
            O => \N__6427\,
            I => \N__6418\
        );

    \I__1405\ : InMux
    port map (
            O => \N__6424\,
            I => \N__6415\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__6421\,
            I => \Instance4.r_CountZ0Z_5\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__6418\,
            I => \Instance4.r_CountZ0Z_5\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__6415\,
            I => \Instance4.r_CountZ0Z_5\
        );

    \I__1401\ : InMux
    port map (
            O => \N__6408\,
            I => \N__6405\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__6405\,
            I => \Instance4.r_Count13_7\
        );

    \I__1399\ : CascadeMux
    port map (
            O => \N__6402\,
            I => \Instance4.r_Count13_13_cascade_\
        );

    \I__1398\ : InMux
    port map (
            O => \N__6399\,
            I => \N__6396\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__6396\,
            I => \N__6393\
        );

    \I__1396\ : Odrv4
    port map (
            O => \N__6393\,
            I => \Instance4.r_Count13_12\
        );

    \I__1395\ : CascadeMux
    port map (
            O => \N__6390\,
            I => \N__6385\
        );

    \I__1394\ : InMux
    port map (
            O => \N__6389\,
            I => \N__6382\
        );

    \I__1393\ : InMux
    port map (
            O => \N__6388\,
            I => \N__6377\
        );

    \I__1392\ : InMux
    port map (
            O => \N__6385\,
            I => \N__6377\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__6382\,
            I => \Instance4.r_CountZ0Z_14\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__6377\,
            I => \Instance4.r_CountZ0Z_14\
        );

    \I__1389\ : InMux
    port map (
            O => \N__6372\,
            I => \N__6367\
        );

    \I__1388\ : InMux
    port map (
            O => \N__6371\,
            I => \N__6362\
        );

    \I__1387\ : InMux
    port map (
            O => \N__6370\,
            I => \N__6362\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__6367\,
            I => \Instance4.r_CountZ0Z_17\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__6362\,
            I => \Instance4.r_CountZ0Z_17\
        );

    \I__1384\ : InMux
    port map (
            O => \N__6357\,
            I => \N__6354\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__6354\,
            I => \Instance4.r_Count13_4\
        );

    \I__1382\ : InMux
    port map (
            O => \N__6351\,
            I => \N__6346\
        );

    \I__1381\ : InMux
    port map (
            O => \N__6350\,
            I => \N__6341\
        );

    \I__1380\ : InMux
    port map (
            O => \N__6349\,
            I => \N__6341\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__6346\,
            I => \Instance4.r_CountZ0Z_11\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__6341\,
            I => \Instance4.r_CountZ0Z_11\
        );

    \I__1377\ : CascadeMux
    port map (
            O => \N__6336\,
            I => \N__6331\
        );

    \I__1376\ : InMux
    port map (
            O => \N__6335\,
            I => \N__6328\
        );

    \I__1375\ : InMux
    port map (
            O => \N__6334\,
            I => \N__6323\
        );

    \I__1374\ : InMux
    port map (
            O => \N__6331\,
            I => \N__6323\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__6328\,
            I => \Instance4.r_CountZ0Z_10\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__6323\,
            I => \Instance4.r_CountZ0Z_10\
        );

    \I__1371\ : InMux
    port map (
            O => \N__6318\,
            I => \N__6313\
        );

    \I__1370\ : InMux
    port map (
            O => \N__6317\,
            I => \N__6310\
        );

    \I__1369\ : InMux
    port map (
            O => \N__6316\,
            I => \N__6307\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__6313\,
            I => \Instance4.r_CountZ0Z_9\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__6310\,
            I => \Instance4.r_CountZ0Z_9\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__6307\,
            I => \Instance4.r_CountZ0Z_9\
        );

    \I__1365\ : InMux
    port map (
            O => \N__6300\,
            I => \N__6295\
        );

    \I__1364\ : InMux
    port map (
            O => \N__6299\,
            I => \N__6292\
        );

    \I__1363\ : InMux
    port map (
            O => \N__6298\,
            I => \N__6289\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__6295\,
            I => \Instance4.r_CountZ0Z_13\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__6292\,
            I => \Instance4.r_CountZ0Z_13\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__6289\,
            I => \Instance4.r_CountZ0Z_13\
        );

    \I__1359\ : InMux
    port map (
            O => \N__6282\,
            I => \N__6277\
        );

    \I__1358\ : InMux
    port map (
            O => \N__6281\,
            I => \N__6274\
        );

    \I__1357\ : InMux
    port map (
            O => \N__6280\,
            I => \N__6271\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__6277\,
            I => \Instance4.r_CountZ0Z_12\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__6274\,
            I => \Instance4.r_CountZ0Z_12\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__6271\,
            I => \Instance4.r_CountZ0Z_12\
        );

    \I__1353\ : CascadeMux
    port map (
            O => \N__6264\,
            I => \Instance4.un1_r_Count_10lto11_1_cascade_\
        );

    \I__1352\ : InMux
    port map (
            O => \N__6261\,
            I => \N__6258\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__6258\,
            I => \Instance4.un1_r_Count_10lt11_0\
        );

    \I__1350\ : InMux
    port map (
            O => \N__6255\,
            I => \N__6249\
        );

    \I__1349\ : InMux
    port map (
            O => \N__6254\,
            I => \N__6249\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__6249\,
            I => \N__6246\
        );

    \I__1347\ : Span4Mux_v
    port map (
            O => \N__6246\,
            I => \N__6243\
        );

    \I__1346\ : Span4Mux_h
    port map (
            O => \N__6243\,
            I => \N__6240\
        );

    \I__1345\ : Odrv4
    port map (
            O => \N__6240\,
            I => \i_Switch_4_c\
        );

    \I__1344\ : InMux
    port map (
            O => \N__6237\,
            I => \N__6231\
        );

    \I__1343\ : InMux
    port map (
            O => \N__6236\,
            I => \N__6231\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__6231\,
            I => \N__6228\
        );

    \I__1341\ : Span4Mux_v
    port map (
            O => \N__6228\,
            I => \N__6223\
        );

    \I__1340\ : InMux
    port map (
            O => \N__6227\,
            I => \N__6218\
        );

    \I__1339\ : InMux
    port map (
            O => \N__6226\,
            I => \N__6218\
        );

    \I__1338\ : Odrv4
    port map (
            O => \N__6223\,
            I => \w_Switch_4\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__6218\,
            I => \w_Switch_4\
        );

    \I__1336\ : CascadeMux
    port map (
            O => \N__6213\,
            I => \Instance4.un1_r_Count_10lt17_cascade_\
        );

    \I__1335\ : InMux
    port map (
            O => \N__6210\,
            I => \N__6207\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__6207\,
            I => \Instance4.un1_r_Count_10lto17_1\
        );

    \I__1333\ : IoInMux
    port map (
            O => \N__6204\,
            I => \N__6201\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__6201\,
            I => \N__6198\
        );

    \I__1331\ : Span12Mux_s1_v
    port map (
            O => \N__6198\,
            I => \N__6195\
        );

    \I__1330\ : Odrv12
    port map (
            O => \N__6195\,
            I => \Instance4.r_Count12_i\
        );

    \I__1329\ : InMux
    port map (
            O => \N__6192\,
            I => \bfn_6_12_0_\
        );

    \I__1328\ : InMux
    port map (
            O => \N__6189\,
            I => \N__6184\
        );

    \I__1327\ : InMux
    port map (
            O => \N__6188\,
            I => \N__6181\
        );

    \I__1326\ : InMux
    port map (
            O => \N__6187\,
            I => \N__6178\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__6184\,
            I => \Instance2.r_CountZ0Z_17\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__6181\,
            I => \Instance2.r_CountZ0Z_17\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__6178\,
            I => \Instance2.r_CountZ0Z_17\
        );

    \I__1322\ : CascadeMux
    port map (
            O => \N__6171\,
            I => \N__6167\
        );

    \I__1321\ : InMux
    port map (
            O => \N__6170\,
            I => \N__6162\
        );

    \I__1320\ : InMux
    port map (
            O => \N__6167\,
            I => \N__6159\
        );

    \I__1319\ : InMux
    port map (
            O => \N__6166\,
            I => \N__6154\
        );

    \I__1318\ : InMux
    port map (
            O => \N__6165\,
            I => \N__6154\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__6162\,
            I => \N__6149\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__6159\,
            I => \N__6149\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__6154\,
            I => \Instance2.r_Count_0_0\
        );

    \I__1314\ : Odrv4
    port map (
            O => \N__6149\,
            I => \Instance2.r_Count_0_0\
        );

    \I__1313\ : InMux
    port map (
            O => \N__6144\,
            I => \N__6139\
        );

    \I__1312\ : CascadeMux
    port map (
            O => \N__6143\,
            I => \N__6136\
        );

    \I__1311\ : InMux
    port map (
            O => \N__6142\,
            I => \N__6133\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__6139\,
            I => \N__6130\
        );

    \I__1309\ : InMux
    port map (
            O => \N__6136\,
            I => \N__6127\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__6133\,
            I => \Instance2.r_Count_0_1\
        );

    \I__1307\ : Odrv4
    port map (
            O => \N__6130\,
            I => \Instance2.r_Count_0_1\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__6127\,
            I => \Instance2.r_Count_0_1\
        );

    \I__1305\ : SRMux
    port map (
            O => \N__6120\,
            I => \N__6111\
        );

    \I__1304\ : SRMux
    port map (
            O => \N__6119\,
            I => \N__6111\
        );

    \I__1303\ : SRMux
    port map (
            O => \N__6118\,
            I => \N__6111\
        );

    \I__1302\ : GlobalMux
    port map (
            O => \N__6111\,
            I => \N__6108\
        );

    \I__1301\ : gio2CtrlBuf
    port map (
            O => \N__6108\,
            I => \Instance2.r_Count12_i_g\
        );

    \I__1300\ : InMux
    port map (
            O => \N__6105\,
            I => \N__6102\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__6102\,
            I => \N__6099\
        );

    \I__1298\ : Span4Mux_v
    port map (
            O => \N__6099\,
            I => \N__6095\
        );

    \I__1297\ : InMux
    port map (
            O => \N__6098\,
            I => \N__6092\
        );

    \I__1296\ : Odrv4
    port map (
            O => \N__6095\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__6092\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1294\ : IoInMux
    port map (
            O => \N__6087\,
            I => \N__6084\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__6084\,
            I => \N__6081\
        );

    \I__1292\ : Odrv12
    port map (
            O => \N__6081\,
            I => \r_HexEncode_i_0_3\
        );

    \I__1291\ : InMux
    port map (
            O => \N__6078\,
            I => \N__6073\
        );

    \I__1290\ : InMux
    port map (
            O => \N__6077\,
            I => \N__6068\
        );

    \I__1289\ : InMux
    port map (
            O => \N__6076\,
            I => \N__6068\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__6073\,
            I => \N__6061\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__6068\,
            I => \N__6061\
        );

    \I__1286\ : InMux
    port map (
            O => \N__6067\,
            I => \N__6054\
        );

    \I__1285\ : InMux
    port map (
            O => \N__6066\,
            I => \N__6054\
        );

    \I__1284\ : Span4Mux_h
    port map (
            O => \N__6061\,
            I => \N__6051\
        );

    \I__1283\ : InMux
    port map (
            O => \N__6060\,
            I => \N__6046\
        );

    \I__1282\ : InMux
    port map (
            O => \N__6059\,
            I => \N__6046\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__6054\,
            I => \N__6043\
        );

    \I__1280\ : Span4Mux_h
    port map (
            O => \N__6051\,
            I => \N__6040\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__6046\,
            I => \sevseglZ0Z_2\
        );

    \I__1278\ : Odrv4
    port map (
            O => \N__6043\,
            I => \sevseglZ0Z_2\
        );

    \I__1277\ : Odrv4
    port map (
            O => \N__6040\,
            I => \sevseglZ0Z_2\
        );

    \I__1276\ : InMux
    port map (
            O => \N__6033\,
            I => \N__6025\
        );

    \I__1275\ : InMux
    port map (
            O => \N__6032\,
            I => \N__6025\
        );

    \I__1274\ : InMux
    port map (
            O => \N__6031\,
            I => \N__6022\
        );

    \I__1273\ : CascadeMux
    port map (
            O => \N__6030\,
            I => \N__6019\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__6025\,
            I => \N__6011\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__6022\,
            I => \N__6011\
        );

    \I__1270\ : InMux
    port map (
            O => \N__6019\,
            I => \N__6006\
        );

    \I__1269\ : InMux
    port map (
            O => \N__6018\,
            I => \N__6006\
        );

    \I__1268\ : InMux
    port map (
            O => \N__6017\,
            I => \N__6001\
        );

    \I__1267\ : InMux
    port map (
            O => \N__6016\,
            I => \N__6001\
        );

    \I__1266\ : Span4Mux_s3_v
    port map (
            O => \N__6011\,
            I => \N__5998\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__6006\,
            I => \sevseglZ0Z_1\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__6001\,
            I => \sevseglZ0Z_1\
        );

    \I__1263\ : Odrv4
    port map (
            O => \N__5998\,
            I => \sevseglZ0Z_1\
        );

    \I__1262\ : CascadeMux
    port map (
            O => \N__5991\,
            I => \N__5986\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__5990\,
            I => \N__5983\
        );

    \I__1260\ : CascadeMux
    port map (
            O => \N__5989\,
            I => \N__5980\
        );

    \I__1259\ : InMux
    port map (
            O => \N__5986\,
            I => \N__5975\
        );

    \I__1258\ : InMux
    port map (
            O => \N__5983\,
            I => \N__5975\
        );

    \I__1257\ : InMux
    port map (
            O => \N__5980\,
            I => \N__5972\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__5975\,
            I => \N__5964\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__5972\,
            I => \N__5964\
        );

    \I__1254\ : CascadeMux
    port map (
            O => \N__5971\,
            I => \N__5960\
        );

    \I__1253\ : CascadeMux
    port map (
            O => \N__5970\,
            I => \N__5957\
        );

    \I__1252\ : CascadeMux
    port map (
            O => \N__5969\,
            I => \N__5954\
        );

    \I__1251\ : Span4Mux_h
    port map (
            O => \N__5964\,
            I => \N__5951\
        );

    \I__1250\ : InMux
    port map (
            O => \N__5963\,
            I => \N__5946\
        );

    \I__1249\ : InMux
    port map (
            O => \N__5960\,
            I => \N__5946\
        );

    \I__1248\ : InMux
    port map (
            O => \N__5957\,
            I => \N__5941\
        );

    \I__1247\ : InMux
    port map (
            O => \N__5954\,
            I => \N__5941\
        );

    \I__1246\ : Odrv4
    port map (
            O => \N__5951\,
            I => \sevseglZ0Z_3\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__5946\,
            I => \sevseglZ0Z_3\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__5941\,
            I => \sevseglZ0Z_3\
        );

    \I__1243\ : InMux
    port map (
            O => \N__5934\,
            I => \N__5928\
        );

    \I__1242\ : InMux
    port map (
            O => \N__5933\,
            I => \N__5928\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__5928\,
            I => \N__5924\
        );

    \I__1240\ : InMux
    port map (
            O => \N__5927\,
            I => \N__5921\
        );

    \I__1239\ : Span4Mux_h
    port map (
            O => \N__5924\,
            I => \N__5916\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__5921\,
            I => \N__5916\
        );

    \I__1237\ : Span4Mux_h
    port map (
            O => \N__5916\,
            I => \N__5909\
        );

    \I__1236\ : InMux
    port map (
            O => \N__5915\,
            I => \N__5904\
        );

    \I__1235\ : InMux
    port map (
            O => \N__5914\,
            I => \N__5904\
        );

    \I__1234\ : InMux
    port map (
            O => \N__5913\,
            I => \N__5899\
        );

    \I__1233\ : InMux
    port map (
            O => \N__5912\,
            I => \N__5899\
        );

    \I__1232\ : Odrv4
    port map (
            O => \N__5909\,
            I => \sevseglZ0Z_0\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__5904\,
            I => \sevseglZ0Z_0\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__5899\,
            I => \sevseglZ0Z_0\
        );

    \I__1229\ : IoInMux
    port map (
            O => \N__5892\,
            I => \N__5889\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__5889\,
            I => \N__5886\
        );

    \I__1227\ : Odrv4
    port map (
            O => \N__5886\,
            I => \r_HexEncode_i_0_2\
        );

    \I__1226\ : InMux
    port map (
            O => \N__5883\,
            I => \N__5878\
        );

    \I__1225\ : InMux
    port map (
            O => \N__5882\,
            I => \N__5875\
        );

    \I__1224\ : InMux
    port map (
            O => \N__5881\,
            I => \N__5872\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__5878\,
            I => \Instance4.r_CountZ0Z_1\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__5875\,
            I => \Instance4.r_CountZ0Z_1\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__5872\,
            I => \Instance4.r_CountZ0Z_1\
        );

    \I__1220\ : InMux
    port map (
            O => \N__5865\,
            I => \N__5861\
        );

    \I__1219\ : InMux
    port map (
            O => \N__5864\,
            I => \N__5858\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__5861\,
            I => \Instance4.r_CountZ0Z_2\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__5858\,
            I => \Instance4.r_CountZ0Z_2\
        );

    \I__1216\ : CascadeMux
    port map (
            O => \N__5853\,
            I => \N__5849\
        );

    \I__1215\ : InMux
    port map (
            O => \N__5852\,
            I => \N__5846\
        );

    \I__1214\ : InMux
    port map (
            O => \N__5849\,
            I => \N__5843\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__5846\,
            I => \Instance4.r_CountZ0Z_3\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__5843\,
            I => \Instance4.r_CountZ0Z_3\
        );

    \I__1211\ : InMux
    port map (
            O => \N__5838\,
            I => \N__5833\
        );

    \I__1210\ : InMux
    port map (
            O => \N__5837\,
            I => \N__5828\
        );

    \I__1209\ : InMux
    port map (
            O => \N__5836\,
            I => \N__5828\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__5833\,
            I => \Instance4.r_CountZ0Z_4\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__5828\,
            I => \Instance4.r_CountZ0Z_4\
        );

    \I__1206\ : CascadeMux
    port map (
            O => \N__5823\,
            I => \N__5820\
        );

    \I__1205\ : InMux
    port map (
            O => \N__5820\,
            I => \N__5815\
        );

    \I__1204\ : InMux
    port map (
            O => \N__5819\,
            I => \N__5812\
        );

    \I__1203\ : InMux
    port map (
            O => \N__5818\,
            I => \N__5809\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__5815\,
            I => \Instance4.r_CountZ0Z_7\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__5812\,
            I => \Instance4.r_CountZ0Z_7\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__5809\,
            I => \Instance4.r_CountZ0Z_7\
        );

    \I__1199\ : InMux
    port map (
            O => \N__5802\,
            I => \N__5797\
        );

    \I__1198\ : InMux
    port map (
            O => \N__5801\,
            I => \N__5792\
        );

    \I__1197\ : InMux
    port map (
            O => \N__5800\,
            I => \N__5792\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__5797\,
            I => \Instance2.r_CountZ0Z_9\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__5792\,
            I => \Instance2.r_CountZ0Z_9\
        );

    \I__1194\ : InMux
    port map (
            O => \N__5787\,
            I => \bfn_6_11_0_\
        );

    \I__1193\ : InMux
    port map (
            O => \N__5784\,
            I => \N__5779\
        );

    \I__1192\ : InMux
    port map (
            O => \N__5783\,
            I => \N__5776\
        );

    \I__1191\ : InMux
    port map (
            O => \N__5782\,
            I => \N__5773\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__5779\,
            I => \N__5770\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__5776\,
            I => \Instance2.r_CountZ0Z_10\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__5773\,
            I => \Instance2.r_CountZ0Z_10\
        );

    \I__1187\ : Odrv4
    port map (
            O => \N__5770\,
            I => \Instance2.r_CountZ0Z_10\
        );

    \I__1186\ : InMux
    port map (
            O => \N__5763\,
            I => \Instance2.r_Count_2_cry_9\
        );

    \I__1185\ : CascadeMux
    port map (
            O => \N__5760\,
            I => \N__5755\
        );

    \I__1184\ : InMux
    port map (
            O => \N__5759\,
            I => \N__5752\
        );

    \I__1183\ : InMux
    port map (
            O => \N__5758\,
            I => \N__5749\
        );

    \I__1182\ : InMux
    port map (
            O => \N__5755\,
            I => \N__5746\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__5752\,
            I => \Instance2.r_CountZ0Z_11\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__5749\,
            I => \Instance2.r_CountZ0Z_11\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__5746\,
            I => \Instance2.r_CountZ0Z_11\
        );

    \I__1178\ : InMux
    port map (
            O => \N__5739\,
            I => \Instance2.r_Count_2_cry_10\
        );

    \I__1177\ : InMux
    port map (
            O => \N__5736\,
            I => \N__5731\
        );

    \I__1176\ : InMux
    port map (
            O => \N__5735\,
            I => \N__5728\
        );

    \I__1175\ : InMux
    port map (
            O => \N__5734\,
            I => \N__5725\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__5731\,
            I => \Instance2.r_CountZ0Z_12\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__5728\,
            I => \Instance2.r_CountZ0Z_12\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__5725\,
            I => \Instance2.r_CountZ0Z_12\
        );

    \I__1171\ : InMux
    port map (
            O => \N__5718\,
            I => \Instance2.r_Count_2_cry_11\
        );

    \I__1170\ : CascadeMux
    port map (
            O => \N__5715\,
            I => \N__5711\
        );

    \I__1169\ : InMux
    port map (
            O => \N__5714\,
            I => \N__5707\
        );

    \I__1168\ : InMux
    port map (
            O => \N__5711\,
            I => \N__5702\
        );

    \I__1167\ : InMux
    port map (
            O => \N__5710\,
            I => \N__5702\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__5707\,
            I => \Instance2.r_CountZ0Z_13\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__5702\,
            I => \Instance2.r_CountZ0Z_13\
        );

    \I__1164\ : InMux
    port map (
            O => \N__5697\,
            I => \Instance2.r_Count_2_cry_12\
        );

    \I__1163\ : CascadeMux
    port map (
            O => \N__5694\,
            I => \N__5689\
        );

    \I__1162\ : InMux
    port map (
            O => \N__5693\,
            I => \N__5686\
        );

    \I__1161\ : InMux
    port map (
            O => \N__5692\,
            I => \N__5683\
        );

    \I__1160\ : InMux
    port map (
            O => \N__5689\,
            I => \N__5680\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__5686\,
            I => \Instance2.r_CountZ0Z_14\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__5683\,
            I => \Instance2.r_CountZ0Z_14\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__5680\,
            I => \Instance2.r_CountZ0Z_14\
        );

    \I__1156\ : InMux
    port map (
            O => \N__5673\,
            I => \Instance2.r_Count_2_cry_13\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__5670\,
            I => \N__5666\
        );

    \I__1154\ : InMux
    port map (
            O => \N__5669\,
            I => \N__5662\
        );

    \I__1153\ : InMux
    port map (
            O => \N__5666\,
            I => \N__5659\
        );

    \I__1152\ : InMux
    port map (
            O => \N__5665\,
            I => \N__5656\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__5662\,
            I => \Instance2.r_CountZ0Z_15\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__5659\,
            I => \Instance2.r_CountZ0Z_15\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__5656\,
            I => \Instance2.r_CountZ0Z_15\
        );

    \I__1148\ : InMux
    port map (
            O => \N__5649\,
            I => \Instance2.r_Count_2_cry_14\
        );

    \I__1147\ : InMux
    port map (
            O => \N__5646\,
            I => \N__5642\
        );

    \I__1146\ : InMux
    port map (
            O => \N__5645\,
            I => \N__5638\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__5642\,
            I => \N__5635\
        );

    \I__1144\ : InMux
    port map (
            O => \N__5641\,
            I => \N__5632\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__5638\,
            I => \Instance2.r_CountZ0Z_16\
        );

    \I__1142\ : Odrv4
    port map (
            O => \N__5635\,
            I => \Instance2.r_CountZ0Z_16\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__5632\,
            I => \Instance2.r_CountZ0Z_16\
        );

    \I__1140\ : InMux
    port map (
            O => \N__5625\,
            I => \Instance2.r_Count_2_cry_15\
        );

    \I__1139\ : SRMux
    port map (
            O => \N__5622\,
            I => \N__5610\
        );

    \I__1138\ : SRMux
    port map (
            O => \N__5621\,
            I => \N__5610\
        );

    \I__1137\ : SRMux
    port map (
            O => \N__5620\,
            I => \N__5610\
        );

    \I__1136\ : SRMux
    port map (
            O => \N__5619\,
            I => \N__5610\
        );

    \I__1135\ : GlobalMux
    port map (
            O => \N__5610\,
            I => \N__5607\
        );

    \I__1134\ : gio2CtrlBuf
    port map (
            O => \N__5607\,
            I => \Instance4.r_Count12_i_g\
        );

    \I__1133\ : InMux
    port map (
            O => \N__5604\,
            I => \N__5600\
        );

    \I__1132\ : InMux
    port map (
            O => \N__5603\,
            I => \N__5597\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__5600\,
            I => \Instance2.r_Count_0_2\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__5597\,
            I => \Instance2.r_Count_0_2\
        );

    \I__1129\ : InMux
    port map (
            O => \N__5592\,
            I => \Instance2.r_Count_2_cry_1\
        );

    \I__1128\ : InMux
    port map (
            O => \N__5589\,
            I => \N__5586\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__5586\,
            I => \N__5583\
        );

    \I__1126\ : Span4Mux_h
    port map (
            O => \N__5583\,
            I => \N__5579\
        );

    \I__1125\ : InMux
    port map (
            O => \N__5582\,
            I => \N__5576\
        );

    \I__1124\ : Odrv4
    port map (
            O => \N__5579\,
            I => \Instance2.r_Count_0_3\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__5576\,
            I => \Instance2.r_Count_0_3\
        );

    \I__1122\ : InMux
    port map (
            O => \N__5571\,
            I => \Instance2.r_Count_2_cry_2\
        );

    \I__1121\ : InMux
    port map (
            O => \N__5568\,
            I => \N__5563\
        );

    \I__1120\ : InMux
    port map (
            O => \N__5567\,
            I => \N__5560\
        );

    \I__1119\ : InMux
    port map (
            O => \N__5566\,
            I => \N__5557\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__5563\,
            I => \N__5552\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__5560\,
            I => \N__5552\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__5557\,
            I => \Instance2.r_CountZ0Z_4\
        );

    \I__1115\ : Odrv4
    port map (
            O => \N__5552\,
            I => \Instance2.r_CountZ0Z_4\
        );

    \I__1114\ : InMux
    port map (
            O => \N__5547\,
            I => \Instance2.r_Count_2_cry_3\
        );

    \I__1113\ : InMux
    port map (
            O => \N__5544\,
            I => \N__5539\
        );

    \I__1112\ : InMux
    port map (
            O => \N__5543\,
            I => \N__5534\
        );

    \I__1111\ : InMux
    port map (
            O => \N__5542\,
            I => \N__5534\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__5539\,
            I => \Instance2.r_CountZ0Z_5\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__5534\,
            I => \Instance2.r_CountZ0Z_5\
        );

    \I__1108\ : InMux
    port map (
            O => \N__5529\,
            I => \Instance2.r_Count_2_cry_4\
        );

    \I__1107\ : InMux
    port map (
            O => \N__5526\,
            I => \N__5521\
        );

    \I__1106\ : InMux
    port map (
            O => \N__5525\,
            I => \N__5518\
        );

    \I__1105\ : InMux
    port map (
            O => \N__5524\,
            I => \N__5515\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__5521\,
            I => \Instance2.r_CountZ0Z_6\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__5518\,
            I => \Instance2.r_CountZ0Z_6\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__5515\,
            I => \Instance2.r_CountZ0Z_6\
        );

    \I__1101\ : InMux
    port map (
            O => \N__5508\,
            I => \Instance2.r_Count_2_cry_5\
        );

    \I__1100\ : CascadeMux
    port map (
            O => \N__5505\,
            I => \N__5500\
        );

    \I__1099\ : InMux
    port map (
            O => \N__5504\,
            I => \N__5497\
        );

    \I__1098\ : InMux
    port map (
            O => \N__5503\,
            I => \N__5494\
        );

    \I__1097\ : InMux
    port map (
            O => \N__5500\,
            I => \N__5491\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__5497\,
            I => \Instance2.r_CountZ0Z_7\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__5494\,
            I => \Instance2.r_CountZ0Z_7\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__5491\,
            I => \Instance2.r_CountZ0Z_7\
        );

    \I__1093\ : InMux
    port map (
            O => \N__5484\,
            I => \Instance2.r_Count_2_cry_6\
        );

    \I__1092\ : InMux
    port map (
            O => \N__5481\,
            I => \N__5476\
        );

    \I__1091\ : InMux
    port map (
            O => \N__5480\,
            I => \N__5471\
        );

    \I__1090\ : InMux
    port map (
            O => \N__5479\,
            I => \N__5471\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__5476\,
            I => \Instance2.r_CountZ0Z_8\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__5471\,
            I => \Instance2.r_CountZ0Z_8\
        );

    \I__1087\ : InMux
    port map (
            O => \N__5466\,
            I => \Instance2.r_Count_2_cry_7\
        );

    \I__1086\ : InMux
    port map (
            O => \N__5463\,
            I => \bfn_6_8_0_\
        );

    \I__1085\ : InMux
    port map (
            O => \N__5460\,
            I => \Instance4.r_Count_2_cry_9\
        );

    \I__1084\ : InMux
    port map (
            O => \N__5457\,
            I => \Instance4.r_Count_2_cry_10\
        );

    \I__1083\ : InMux
    port map (
            O => \N__5454\,
            I => \Instance4.r_Count_2_cry_11\
        );

    \I__1082\ : InMux
    port map (
            O => \N__5451\,
            I => \Instance4.r_Count_2_cry_12\
        );

    \I__1081\ : InMux
    port map (
            O => \N__5448\,
            I => \Instance4.r_Count_2_cry_13\
        );

    \I__1080\ : InMux
    port map (
            O => \N__5445\,
            I => \Instance4.r_Count_2_cry_14\
        );

    \I__1079\ : InMux
    port map (
            O => \N__5442\,
            I => \Instance4.r_Count_2_cry_15\
        );

    \I__1078\ : InMux
    port map (
            O => \N__5439\,
            I => \bfn_6_9_0_\
        );

    \I__1077\ : InMux
    port map (
            O => \N__5436\,
            I => \Instance4.r_Count_2_cry_1\
        );

    \I__1076\ : InMux
    port map (
            O => \N__5433\,
            I => \Instance4.r_Count_2_cry_2\
        );

    \I__1075\ : InMux
    port map (
            O => \N__5430\,
            I => \Instance4.r_Count_2_cry_3\
        );

    \I__1074\ : InMux
    port map (
            O => \N__5427\,
            I => \Instance4.r_Count_2_cry_4\
        );

    \I__1073\ : InMux
    port map (
            O => \N__5424\,
            I => \Instance4.r_Count_2_cry_5\
        );

    \I__1072\ : InMux
    port map (
            O => \N__5421\,
            I => \Instance4.r_Count_2_cry_6\
        );

    \I__1071\ : InMux
    port map (
            O => \N__5418\,
            I => \Instance4.r_Count_2_cry_7\
        );

    \I__1070\ : IoInMux
    port map (
            O => \N__5415\,
            I => \N__5412\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__5412\,
            I => \N__5409\
        );

    \I__1068\ : Odrv4
    port map (
            O => \N__5409\,
            I => \r_HexEncode_i_0_4\
        );

    \I__1067\ : CEMux
    port map (
            O => \N__5406\,
            I => \N__5401\
        );

    \I__1066\ : CEMux
    port map (
            O => \N__5405\,
            I => \N__5397\
        );

    \I__1065\ : CEMux
    port map (
            O => \N__5404\,
            I => \N__5394\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__5401\,
            I => \N__5391\
        );

    \I__1063\ : CEMux
    port map (
            O => \N__5400\,
            I => \N__5388\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__5397\,
            I => \N__5383\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__5394\,
            I => \N__5383\
        );

    \I__1060\ : Span4Mux_v
    port map (
            O => \N__5391\,
            I => \N__5380\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__5388\,
            I => \N__5377\
        );

    \I__1058\ : Span4Mux_h
    port map (
            O => \N__5383\,
            I => \N__5374\
        );

    \I__1057\ : Span4Mux_h
    port map (
            O => \N__5380\,
            I => \N__5369\
        );

    \I__1056\ : Span4Mux_h
    port map (
            O => \N__5377\,
            I => \N__5369\
        );

    \I__1055\ : Odrv4
    port map (
            O => \N__5374\,
            I => \alogicunit.N_35\
        );

    \I__1054\ : Odrv4
    port map (
            O => \N__5369\,
            I => \alogicunit.N_35\
        );

    \I__1053\ : InMux
    port map (
            O => \N__5364\,
            I => \N__5358\
        );

    \I__1052\ : InMux
    port map (
            O => \N__5363\,
            I => \N__5358\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__5358\,
            I => \N__5352\
        );

    \I__1050\ : InMux
    port map (
            O => \N__5357\,
            I => \N__5347\
        );

    \I__1049\ : InMux
    port map (
            O => \N__5356\,
            I => \N__5347\
        );

    \I__1048\ : InMux
    port map (
            O => \N__5355\,
            I => \N__5344\
        );

    \I__1047\ : Odrv4
    port map (
            O => \N__5352\,
            I => \alogicunit.result24_iZ0\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__5347\,
            I => \alogicunit.result24_iZ0\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__5344\,
            I => \alogicunit.result24_iZ0\
        );

    \I__1044\ : InMux
    port map (
            O => \N__5337\,
            I => \N__5332\
        );

    \I__1043\ : CascadeMux
    port map (
            O => \N__5336\,
            I => \N__5329\
        );

    \I__1042\ : CascadeMux
    port map (
            O => \N__5335\,
            I => \N__5324\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__5332\,
            I => \N__5316\
        );

    \I__1040\ : InMux
    port map (
            O => \N__5329\,
            I => \N__5312\
        );

    \I__1039\ : InMux
    port map (
            O => \N__5328\,
            I => \N__5307\
        );

    \I__1038\ : InMux
    port map (
            O => \N__5327\,
            I => \N__5307\
        );

    \I__1037\ : InMux
    port map (
            O => \N__5324\,
            I => \N__5304\
        );

    \I__1036\ : CascadeMux
    port map (
            O => \N__5323\,
            I => \N__5298\
        );

    \I__1035\ : InMux
    port map (
            O => \N__5322\,
            I => \N__5291\
        );

    \I__1034\ : InMux
    port map (
            O => \N__5321\,
            I => \N__5284\
        );

    \I__1033\ : InMux
    port map (
            O => \N__5320\,
            I => \N__5284\
        );

    \I__1032\ : InMux
    port map (
            O => \N__5319\,
            I => \N__5284\
        );

    \I__1031\ : Span4Mux_h
    port map (
            O => \N__5316\,
            I => \N__5281\
        );

    \I__1030\ : InMux
    port map (
            O => \N__5315\,
            I => \N__5278\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__5312\,
            I => \N__5271\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__5307\,
            I => \N__5271\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__5304\,
            I => \N__5271\
        );

    \I__1026\ : InMux
    port map (
            O => \N__5303\,
            I => \N__5260\
        );

    \I__1025\ : InMux
    port map (
            O => \N__5302\,
            I => \N__5260\
        );

    \I__1024\ : InMux
    port map (
            O => \N__5301\,
            I => \N__5260\
        );

    \I__1023\ : InMux
    port map (
            O => \N__5298\,
            I => \N__5260\
        );

    \I__1022\ : InMux
    port map (
            O => \N__5297\,
            I => \N__5260\
        );

    \I__1021\ : InMux
    port map (
            O => \N__5296\,
            I => \N__5257\
        );

    \I__1020\ : InMux
    port map (
            O => \N__5295\,
            I => \N__5252\
        );

    \I__1019\ : InMux
    port map (
            O => \N__5294\,
            I => \N__5252\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__5291\,
            I => current_state_0
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__5284\,
            I => current_state_0
        );

    \I__1016\ : Odrv4
    port map (
            O => \N__5281\,
            I => current_state_0
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__5278\,
            I => current_state_0
        );

    \I__1014\ : Odrv4
    port map (
            O => \N__5271\,
            I => current_state_0
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__5260\,
            I => current_state_0
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__5257\,
            I => current_state_0
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__5252\,
            I => current_state_0
        );

    \I__1010\ : CascadeMux
    port map (
            O => \N__5235\,
            I => \N__5231\
        );

    \I__1009\ : CascadeMux
    port map (
            O => \N__5234\,
            I => \N__5228\
        );

    \I__1008\ : InMux
    port map (
            O => \N__5231\,
            I => \N__5217\
        );

    \I__1007\ : InMux
    port map (
            O => \N__5228\,
            I => \N__5217\
        );

    \I__1006\ : InMux
    port map (
            O => \N__5227\,
            I => \N__5214\
        );

    \I__1005\ : InMux
    port map (
            O => \N__5226\,
            I => \N__5211\
        );

    \I__1004\ : CascadeMux
    port map (
            O => \N__5225\,
            I => \N__5203\
        );

    \I__1003\ : CascadeMux
    port map (
            O => \N__5224\,
            I => \N__5197\
        );

    \I__1002\ : InMux
    port map (
            O => \N__5223\,
            I => \N__5194\
        );

    \I__1001\ : InMux
    port map (
            O => \N__5222\,
            I => \N__5191\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__5217\,
            I => \N__5186\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__5214\,
            I => \N__5186\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__5211\,
            I => \N__5183\
        );

    \I__997\ : InMux
    port map (
            O => \N__5210\,
            I => \N__5170\
        );

    \I__996\ : InMux
    port map (
            O => \N__5209\,
            I => \N__5170\
        );

    \I__995\ : InMux
    port map (
            O => \N__5208\,
            I => \N__5170\
        );

    \I__994\ : InMux
    port map (
            O => \N__5207\,
            I => \N__5170\
        );

    \I__993\ : InMux
    port map (
            O => \N__5206\,
            I => \N__5170\
        );

    \I__992\ : InMux
    port map (
            O => \N__5203\,
            I => \N__5170\
        );

    \I__991\ : InMux
    port map (
            O => \N__5202\,
            I => \N__5161\
        );

    \I__990\ : InMux
    port map (
            O => \N__5201\,
            I => \N__5161\
        );

    \I__989\ : InMux
    port map (
            O => \N__5200\,
            I => \N__5161\
        );

    \I__988\ : InMux
    port map (
            O => \N__5197\,
            I => \N__5161\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__5194\,
            I => current_state_1
        );

    \I__986\ : LocalMux
    port map (
            O => \N__5191\,
            I => current_state_1
        );

    \I__985\ : Odrv4
    port map (
            O => \N__5186\,
            I => current_state_1
        );

    \I__984\ : Odrv4
    port map (
            O => \N__5183\,
            I => current_state_1
        );

    \I__983\ : LocalMux
    port map (
            O => \N__5170\,
            I => current_state_1
        );

    \I__982\ : LocalMux
    port map (
            O => \N__5161\,
            I => current_state_1
        );

    \I__981\ : InMux
    port map (
            O => \N__5148\,
            I => \N__5134\
        );

    \I__980\ : InMux
    port map (
            O => \N__5147\,
            I => \N__5134\
        );

    \I__979\ : InMux
    port map (
            O => \N__5146\,
            I => \N__5134\
        );

    \I__978\ : InMux
    port map (
            O => \N__5145\,
            I => \N__5127\
        );

    \I__977\ : InMux
    port map (
            O => \N__5144\,
            I => \N__5122\
        );

    \I__976\ : InMux
    port map (
            O => \N__5143\,
            I => \N__5122\
        );

    \I__975\ : InMux
    port map (
            O => \N__5142\,
            I => \N__5119\
        );

    \I__974\ : CascadeMux
    port map (
            O => \N__5141\,
            I => \N__5115\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__5134\,
            I => \N__5112\
        );

    \I__972\ : CascadeMux
    port map (
            O => \N__5133\,
            I => \N__5108\
        );

    \I__971\ : CascadeMux
    port map (
            O => \N__5132\,
            I => \N__5103\
        );

    \I__970\ : InMux
    port map (
            O => \N__5131\,
            I => \N__5097\
        );

    \I__969\ : InMux
    port map (
            O => \N__5130\,
            I => \N__5094\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__5127\,
            I => \N__5089\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__5122\,
            I => \N__5089\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__5119\,
            I => \N__5086\
        );

    \I__965\ : InMux
    port map (
            O => \N__5118\,
            I => \N__5081\
        );

    \I__964\ : InMux
    port map (
            O => \N__5115\,
            I => \N__5081\
        );

    \I__963\ : Span4Mux_v
    port map (
            O => \N__5112\,
            I => \N__5078\
        );

    \I__962\ : InMux
    port map (
            O => \N__5111\,
            I => \N__5067\
        );

    \I__961\ : InMux
    port map (
            O => \N__5108\,
            I => \N__5067\
        );

    \I__960\ : InMux
    port map (
            O => \N__5107\,
            I => \N__5067\
        );

    \I__959\ : InMux
    port map (
            O => \N__5106\,
            I => \N__5067\
        );

    \I__958\ : InMux
    port map (
            O => \N__5103\,
            I => \N__5067\
        );

    \I__957\ : InMux
    port map (
            O => \N__5102\,
            I => \N__5064\
        );

    \I__956\ : InMux
    port map (
            O => \N__5101\,
            I => \N__5059\
        );

    \I__955\ : InMux
    port map (
            O => \N__5100\,
            I => \N__5059\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__5097\,
            I => current_state_2
        );

    \I__953\ : LocalMux
    port map (
            O => \N__5094\,
            I => current_state_2
        );

    \I__952\ : Odrv4
    port map (
            O => \N__5089\,
            I => current_state_2
        );

    \I__951\ : Odrv4
    port map (
            O => \N__5086\,
            I => current_state_2
        );

    \I__950\ : LocalMux
    port map (
            O => \N__5081\,
            I => current_state_2
        );

    \I__949\ : Odrv4
    port map (
            O => \N__5078\,
            I => current_state_2
        );

    \I__948\ : LocalMux
    port map (
            O => \N__5067\,
            I => current_state_2
        );

    \I__947\ : LocalMux
    port map (
            O => \N__5064\,
            I => current_state_2
        );

    \I__946\ : LocalMux
    port map (
            O => \N__5059\,
            I => current_state_2
        );

    \I__945\ : InMux
    port map (
            O => \N__5040\,
            I => \N__5034\
        );

    \I__944\ : InMux
    port map (
            O => \N__5039\,
            I => \N__5029\
        );

    \I__943\ : InMux
    port map (
            O => \N__5038\,
            I => \N__5029\
        );

    \I__942\ : InMux
    port map (
            O => \N__5037\,
            I => \N__5026\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__5034\,
            I => \N__5013\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__5029\,
            I => \N__5013\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__5026\,
            I => \N__5010\
        );

    \I__938\ : InMux
    port map (
            O => \N__5025\,
            I => \N__5005\
        );

    \I__937\ : InMux
    port map (
            O => \N__5024\,
            I => \N__5005\
        );

    \I__936\ : InMux
    port map (
            O => \N__5023\,
            I => \N__4992\
        );

    \I__935\ : InMux
    port map (
            O => \N__5022\,
            I => \N__4992\
        );

    \I__934\ : InMux
    port map (
            O => \N__5021\,
            I => \N__4992\
        );

    \I__933\ : InMux
    port map (
            O => \N__5020\,
            I => \N__4992\
        );

    \I__932\ : InMux
    port map (
            O => \N__5019\,
            I => \N__4992\
        );

    \I__931\ : InMux
    port map (
            O => \N__5018\,
            I => \N__4992\
        );

    \I__930\ : Span4Mux_v
    port map (
            O => \N__5013\,
            I => \N__4979\
        );

    \I__929\ : Span4Mux_h
    port map (
            O => \N__5010\,
            I => \N__4979\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__5005\,
            I => \N__4979\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__4992\,
            I => \N__4979\
        );

    \I__926\ : InMux
    port map (
            O => \N__4991\,
            I => \N__4970\
        );

    \I__925\ : InMux
    port map (
            O => \N__4990\,
            I => \N__4970\
        );

    \I__924\ : InMux
    port map (
            O => \N__4989\,
            I => \N__4970\
        );

    \I__923\ : InMux
    port map (
            O => \N__4988\,
            I => \N__4970\
        );

    \I__922\ : Odrv4
    port map (
            O => \N__4979\,
            I => current_state_3
        );

    \I__921\ : LocalMux
    port map (
            O => \N__4970\,
            I => current_state_3
        );

    \I__920\ : CEMux
    port map (
            O => \N__4965\,
            I => \N__4960\
        );

    \I__919\ : CascadeMux
    port map (
            O => \N__4964\,
            I => \N__4956\
        );

    \I__918\ : InMux
    port map (
            O => \N__4963\,
            I => \N__4952\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__4960\,
            I => \N__4949\
        );

    \I__916\ : InMux
    port map (
            O => \N__4959\,
            I => \N__4946\
        );

    \I__915\ : InMux
    port map (
            O => \N__4956\,
            I => \N__4941\
        );

    \I__914\ : InMux
    port map (
            O => \N__4955\,
            I => \N__4941\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__4952\,
            I => \N__4938\
        );

    \I__912\ : Span4Mux_s2_v
    port map (
            O => \N__4949\,
            I => \N__4931\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__4946\,
            I => \N__4931\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__4941\,
            I => \N__4931\
        );

    \I__909\ : Odrv4
    port map (
            O => \N__4938\,
            I => \clickZ0Z1\
        );

    \I__908\ : Odrv4
    port map (
            O => \N__4931\,
            I => \clickZ0Z1\
        );

    \I__907\ : InMux
    port map (
            O => \N__4926\,
            I => \N__4923\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__4923\,
            I => \N__4920\
        );

    \I__905\ : Odrv12
    port map (
            O => \N__4920\,
            I => \Instance2.un1_r_Count_10lto17_1\
        );

    \I__904\ : InMux
    port map (
            O => \N__4917\,
            I => \N__4912\
        );

    \I__903\ : InMux
    port map (
            O => \N__4916\,
            I => \N__4909\
        );

    \I__902\ : InMux
    port map (
            O => \N__4915\,
            I => \N__4906\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__4912\,
            I => \N__4903\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__4909\,
            I => \N__4898\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__4906\,
            I => \N__4895\
        );

    \I__898\ : Span12Mux_s4_h
    port map (
            O => \N__4903\,
            I => \N__4892\
        );

    \I__897\ : InMux
    port map (
            O => \N__4902\,
            I => \N__4887\
        );

    \I__896\ : InMux
    port map (
            O => \N__4901\,
            I => \N__4887\
        );

    \I__895\ : Odrv4
    port map (
            O => \N__4898\,
            I => \w_Switch_2\
        );

    \I__894\ : Odrv12
    port map (
            O => \N__4895\,
            I => \w_Switch_2\
        );

    \I__893\ : Odrv12
    port map (
            O => \N__4892\,
            I => \w_Switch_2\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__4887\,
            I => \w_Switch_2\
        );

    \I__891\ : CascadeMux
    port map (
            O => \N__4878\,
            I => \N__4875\
        );

    \I__890\ : InMux
    port map (
            O => \N__4875\,
            I => \N__4872\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__4872\,
            I => \N__4868\
        );

    \I__888\ : InMux
    port map (
            O => \N__4871\,
            I => \N__4865\
        );

    \I__887\ : Span4Mux_s3_v
    port map (
            O => \N__4868\,
            I => \N__4862\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__4865\,
            I => \N__4859\
        );

    \I__885\ : Sp12to4
    port map (
            O => \N__4862\,
            I => \N__4854\
        );

    \I__884\ : Sp12to4
    port map (
            O => \N__4859\,
            I => \N__4854\
        );

    \I__883\ : Span12Mux_v
    port map (
            O => \N__4854\,
            I => \N__4851\
        );

    \I__882\ : Odrv12
    port map (
            O => \N__4851\,
            I => \i_Switch_2_c\
        );

    \I__881\ : InMux
    port map (
            O => \N__4848\,
            I => \N__4845\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__4845\,
            I => \N__4842\
        );

    \I__879\ : Odrv12
    port map (
            O => \N__4842\,
            I => \Instance2.un1_r_Count_10lt17\
        );

    \I__878\ : IoInMux
    port map (
            O => \N__4839\,
            I => \N__4836\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__4836\,
            I => \Instance2.r_Count12_i\
        );

    \I__876\ : InMux
    port map (
            O => \N__4833\,
            I => \N__4830\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__4830\,
            I => \N__4826\
        );

    \I__874\ : InMux
    port map (
            O => \N__4829\,
            I => \N__4823\
        );

    \I__873\ : Odrv12
    port map (
            O => \N__4826\,
            I => \r_SwitchZ0Z_2\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__4823\,
            I => \r_SwitchZ0Z_2\
        );

    \I__871\ : InMux
    port map (
            O => \N__4818\,
            I => \N__4815\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__4815\,
            I => \r_SwitchZ0Z_4\
        );

    \I__869\ : CascadeMux
    port map (
            O => \N__4812\,
            I => \Instance2.click14_sn_cascade_\
        );

    \I__868\ : InMux
    port map (
            O => \N__4809\,
            I => \N__4802\
        );

    \I__867\ : InMux
    port map (
            O => \N__4808\,
            I => \N__4797\
        );

    \I__866\ : InMux
    port map (
            O => \N__4807\,
            I => \N__4797\
        );

    \I__865\ : InMux
    port map (
            O => \N__4806\,
            I => \N__4794\
        );

    \I__864\ : CascadeMux
    port map (
            O => \N__4805\,
            I => \N__4791\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__4802\,
            I => \N__4782\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__4797\,
            I => \N__4782\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__4794\,
            I => \N__4782\
        );

    \I__860\ : InMux
    port map (
            O => \N__4791\,
            I => \N__4774\
        );

    \I__859\ : InMux
    port map (
            O => \N__4790\,
            I => \N__4774\
        );

    \I__858\ : InMux
    port map (
            O => \N__4789\,
            I => \N__4774\
        );

    \I__857\ : Span4Mux_v
    port map (
            O => \N__4782\,
            I => \N__4771\
        );

    \I__856\ : InMux
    port map (
            O => \N__4781\,
            I => \N__4768\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__4774\,
            I => un1_click13_1_sn
        );

    \I__854\ : Odrv4
    port map (
            O => \N__4771\,
            I => un1_click13_1_sn
        );

    \I__853\ : LocalMux
    port map (
            O => \N__4768\,
            I => un1_click13_1_sn
        );

    \I__852\ : InMux
    port map (
            O => \N__4761\,
            I => \N__4757\
        );

    \I__851\ : InMux
    port map (
            O => \N__4760\,
            I => \N__4754\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__4757\,
            I => \N__4751\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__4754\,
            I => \Instance2_un1_click13_3_1\
        );

    \I__848\ : Odrv12
    port map (
            O => \N__4751\,
            I => \Instance2_un1_click13_3_1\
        );

    \I__847\ : InMux
    port map (
            O => \N__4746\,
            I => \N__4743\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__4743\,
            I => \alogicunit.result_RNO_0Z0Z_4\
        );

    \I__845\ : CascadeMux
    port map (
            O => \N__4740\,
            I => \N__4737\
        );

    \I__844\ : InMux
    port map (
            O => \N__4737\,
            I => \N__4734\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__4734\,
            I => \N__4731\
        );

    \I__842\ : Span4Mux_s2_h
    port map (
            O => \N__4731\,
            I => \N__4728\
        );

    \I__841\ : Odrv4
    port map (
            O => \N__4728\,
            I => left_0
        );

    \I__840\ : InMux
    port map (
            O => \N__4725\,
            I => \N__4719\
        );

    \I__839\ : InMux
    port map (
            O => \N__4724\,
            I => \N__4719\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__4719\,
            I => \alogicunit.N_50\
        );

    \I__837\ : InMux
    port map (
            O => \N__4716\,
            I => \N__4713\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__4713\,
            I => \alogicunit.result_RNO_0Z0Z_6\
        );

    \I__835\ : InMux
    port map (
            O => \N__4710\,
            I => \N__4707\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__4707\,
            I => \N__4704\
        );

    \I__833\ : Span4Mux_s2_h
    port map (
            O => \N__4704\,
            I => \N__4701\
        );

    \I__832\ : Odrv4
    port map (
            O => \N__4701\,
            I => left_2
        );

    \I__831\ : InMux
    port map (
            O => \N__4698\,
            I => \N__4694\
        );

    \I__830\ : InMux
    port map (
            O => \N__4697\,
            I => \N__4691\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__4694\,
            I => \alogicunit.un1_a_1_cry_1_c_invZ0\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__4691\,
            I => \alogicunit.un1_a_1_cry_1_c_invZ0\
        );

    \I__827\ : InMux
    port map (
            O => \N__4686\,
            I => \N__4680\
        );

    \I__826\ : InMux
    port map (
            O => \N__4685\,
            I => \N__4680\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__4680\,
            I => \alogicunit.N_102\
        );

    \I__824\ : InMux
    port map (
            O => \N__4677\,
            I => \N__4674\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__4674\,
            I => \Instance2.r_Count13_12\
        );

    \I__822\ : CascadeMux
    port map (
            O => \N__4671\,
            I => \Instance2.r_Count13_13_cascade_\
        );

    \I__821\ : InMux
    port map (
            O => \N__4668\,
            I => \N__4665\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__4665\,
            I => \Instance2.un1_r_Count_10lto11_1\
        );

    \I__819\ : CascadeMux
    port map (
            O => \N__4662\,
            I => \N__4659\
        );

    \I__818\ : InMux
    port map (
            O => \N__4659\,
            I => \N__4656\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__4656\,
            I => \Instance2.r_Count13_10\
        );

    \I__816\ : InMux
    port map (
            O => \N__4653\,
            I => \N__4650\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__4650\,
            I => \Instance2.r_Count13_7\
        );

    \I__814\ : CascadeMux
    port map (
            O => \N__4647\,
            I => \N__4644\
        );

    \I__813\ : InMux
    port map (
            O => \N__4644\,
            I => \N__4638\
        );

    \I__812\ : InMux
    port map (
            O => \N__4643\,
            I => \N__4638\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__4638\,
            I => \alogicunit.N_90\
        );

    \I__810\ : InMux
    port map (
            O => \N__4635\,
            I => \N__4632\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__4632\,
            I => \Instance2.r_Count13_4\
        );

    \I__808\ : CEMux
    port map (
            O => \N__4629\,
            I => \N__4626\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__4626\,
            I => \N__4617\
        );

    \I__806\ : InMux
    port map (
            O => \N__4625\,
            I => \N__4614\
        );

    \I__805\ : InMux
    port map (
            O => \N__4624\,
            I => \N__4607\
        );

    \I__804\ : InMux
    port map (
            O => \N__4623\,
            I => \N__4607\
        );

    \I__803\ : InMux
    port map (
            O => \N__4622\,
            I => \N__4607\
        );

    \I__802\ : InMux
    port map (
            O => \N__4621\,
            I => \N__4599\
        );

    \I__801\ : InMux
    port map (
            O => \N__4620\,
            I => \N__4599\
        );

    \I__800\ : Span4Mux_h
    port map (
            O => \N__4617\,
            I => \N__4594\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__4614\,
            I => \N__4594\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__4607\,
            I => \N__4591\
        );

    \I__797\ : InMux
    port map (
            O => \N__4606\,
            I => \N__4588\
        );

    \I__796\ : InMux
    port map (
            O => \N__4605\,
            I => \N__4583\
        );

    \I__795\ : InMux
    port map (
            O => \N__4604\,
            I => \N__4583\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__4599\,
            I => \N__4575\
        );

    \I__793\ : Span4Mux_v
    port map (
            O => \N__4594\,
            I => \N__4570\
        );

    \I__792\ : Span4Mux_v
    port map (
            O => \N__4591\,
            I => \N__4570\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__4588\,
            I => \N__4567\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__4583\,
            I => \N__4564\
        );

    \I__789\ : InMux
    port map (
            O => \N__4582\,
            I => \N__4557\
        );

    \I__788\ : InMux
    port map (
            O => \N__4581\,
            I => \N__4557\
        );

    \I__787\ : InMux
    port map (
            O => \N__4580\,
            I => \N__4557\
        );

    \I__786\ : InMux
    port map (
            O => \N__4579\,
            I => \N__4552\
        );

    \I__785\ : InMux
    port map (
            O => \N__4578\,
            I => \N__4552\
        );

    \I__784\ : Odrv4
    port map (
            O => \N__4575\,
            I => click13
        );

    \I__783\ : Odrv4
    port map (
            O => \N__4570\,
            I => click13
        );

    \I__782\ : Odrv12
    port map (
            O => \N__4567\,
            I => click13
        );

    \I__781\ : Odrv4
    port map (
            O => \N__4564\,
            I => click13
        );

    \I__780\ : LocalMux
    port map (
            O => \N__4557\,
            I => click13
        );

    \I__779\ : LocalMux
    port map (
            O => \N__4552\,
            I => click13
        );

    \I__778\ : InMux
    port map (
            O => \N__4539\,
            I => \N__4535\
        );

    \I__777\ : InMux
    port map (
            O => \N__4538\,
            I => \N__4532\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__4535\,
            I => \alogicunit.N_49\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__4532\,
            I => \alogicunit.N_49\
        );

    \I__774\ : InMux
    port map (
            O => \N__4527\,
            I => \N__4524\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__4524\,
            I => \N__4521\
        );

    \I__772\ : Span4Mux_s3_h
    port map (
            O => \N__4521\,
            I => \N__4517\
        );

    \I__771\ : InMux
    port map (
            O => \N__4520\,
            I => \N__4514\
        );

    \I__770\ : Odrv4
    port map (
            O => \N__4517\,
            I => \N_28\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__4514\,
            I => \N_28\
        );

    \I__768\ : InMux
    port map (
            O => \N__4509\,
            I => \N__4503\
        );

    \I__767\ : InMux
    port map (
            O => \N__4508\,
            I => \N__4503\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__4503\,
            I => \N__4500\
        );

    \I__765\ : Span4Mux_s3_h
    port map (
            O => \N__4500\,
            I => \N__4497\
        );

    \I__764\ : Odrv4
    port map (
            O => \N__4497\,
            I => \alogicunit.N_41\
        );

    \I__763\ : CascadeMux
    port map (
            O => \N__4494\,
            I => \alogicunit.N_41_cascade_\
        );

    \I__762\ : CascadeMux
    port map (
            O => \N__4491\,
            I => \N__4487\
        );

    \I__761\ : CascadeMux
    port map (
            O => \N__4490\,
            I => \N__4484\
        );

    \I__760\ : InMux
    port map (
            O => \N__4487\,
            I => \N__4481\
        );

    \I__759\ : InMux
    port map (
            O => \N__4484\,
            I => \N__4478\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__4481\,
            I => \N__4475\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__4478\,
            I => \N__4472\
        );

    \I__756\ : Span4Mux_s3_h
    port map (
            O => \N__4475\,
            I => \N__4469\
        );

    \I__755\ : Span4Mux_v
    port map (
            O => \N__4472\,
            I => \N__4466\
        );

    \I__754\ : Odrv4
    port map (
            O => \N__4469\,
            I => \track_RNI9MAL_0_1\
        );

    \I__753\ : Odrv4
    port map (
            O => \N__4466\,
            I => \track_RNI9MAL_0_1\
        );

    \I__752\ : CascadeMux
    port map (
            O => \N__4461\,
            I => \N__4456\
        );

    \I__751\ : InMux
    port map (
            O => \N__4460\,
            I => \N__4450\
        );

    \I__750\ : InMux
    port map (
            O => \N__4459\,
            I => \N__4447\
        );

    \I__749\ : InMux
    port map (
            O => \N__4456\,
            I => \N__4442\
        );

    \I__748\ : InMux
    port map (
            O => \N__4455\,
            I => \N__4442\
        );

    \I__747\ : InMux
    port map (
            O => \N__4454\,
            I => \N__4439\
        );

    \I__746\ : InMux
    port map (
            O => \N__4453\,
            I => \N__4435\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__4450\,
            I => \N__4432\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__4447\,
            I => \N__4429\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__4442\,
            I => \N__4426\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__4439\,
            I => \N__4423\
        );

    \I__741\ : CascadeMux
    port map (
            O => \N__4438\,
            I => \N__4420\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__4435\,
            I => \N__4415\
        );

    \I__739\ : Span4Mux_v
    port map (
            O => \N__4432\,
            I => \N__4410\
        );

    \I__738\ : Span4Mux_v
    port map (
            O => \N__4429\,
            I => \N__4410\
        );

    \I__737\ : Span4Mux_h
    port map (
            O => \N__4426\,
            I => \N__4405\
        );

    \I__736\ : Span4Mux_s3_h
    port map (
            O => \N__4423\,
            I => \N__4405\
        );

    \I__735\ : InMux
    port map (
            O => \N__4420\,
            I => \N__4398\
        );

    \I__734\ : InMux
    port map (
            O => \N__4419\,
            I => \N__4398\
        );

    \I__733\ : InMux
    port map (
            O => \N__4418\,
            I => \N__4398\
        );

    \I__732\ : Odrv12
    port map (
            O => \N__4415\,
            I => \r_CountZ0Z_1\
        );

    \I__731\ : Odrv4
    port map (
            O => \N__4410\,
            I => \r_CountZ0Z_1\
        );

    \I__730\ : Odrv4
    port map (
            O => \N__4405\,
            I => \r_CountZ0Z_1\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__4398\,
            I => \r_CountZ0Z_1\
        );

    \I__728\ : InMux
    port map (
            O => \N__4389\,
            I => \N__4377\
        );

    \I__727\ : InMux
    port map (
            O => \N__4388\,
            I => \N__4377\
        );

    \I__726\ : InMux
    port map (
            O => \N__4387\,
            I => \N__4377\
        );

    \I__725\ : InMux
    port map (
            O => \N__4386\,
            I => \N__4372\
        );

    \I__724\ : InMux
    port map (
            O => \N__4385\,
            I => \N__4372\
        );

    \I__723\ : InMux
    port map (
            O => \N__4384\,
            I => \N__4369\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__4377\,
            I => \N__4366\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__4372\,
            I => \N__4363\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__4369\,
            I => \N__4356\
        );

    \I__719\ : Span4Mux_s3_h
    port map (
            O => \N__4366\,
            I => \N__4353\
        );

    \I__718\ : Span4Mux_s3_h
    port map (
            O => \N__4363\,
            I => \N__4350\
        );

    \I__717\ : InMux
    port map (
            O => \N__4362\,
            I => \N__4341\
        );

    \I__716\ : InMux
    port map (
            O => \N__4361\,
            I => \N__4341\
        );

    \I__715\ : InMux
    port map (
            O => \N__4360\,
            I => \N__4341\
        );

    \I__714\ : InMux
    port map (
            O => \N__4359\,
            I => \N__4341\
        );

    \I__713\ : Odrv12
    port map (
            O => \N__4356\,
            I => \r_CountZ0Z_0\
        );

    \I__712\ : Odrv4
    port map (
            O => \N__4353\,
            I => \r_CountZ0Z_0\
        );

    \I__711\ : Odrv4
    port map (
            O => \N__4350\,
            I => \r_CountZ0Z_0\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__4341\,
            I => \r_CountZ0Z_0\
        );

    \I__709\ : InMux
    port map (
            O => \N__4332\,
            I => \N__4328\
        );

    \I__708\ : InMux
    port map (
            O => \N__4331\,
            I => \N__4324\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__4328\,
            I => \N__4318\
        );

    \I__706\ : InMux
    port map (
            O => \N__4327\,
            I => \N__4315\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__4324\,
            I => \N__4312\
        );

    \I__704\ : InMux
    port map (
            O => \N__4323\,
            I => \N__4307\
        );

    \I__703\ : InMux
    port map (
            O => \N__4322\,
            I => \N__4307\
        );

    \I__702\ : InMux
    port map (
            O => \N__4321\,
            I => \N__4304\
        );

    \I__701\ : Span4Mux_h
    port map (
            O => \N__4318\,
            I => \N__4301\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__4315\,
            I => \N__4298\
        );

    \I__699\ : Span4Mux_s3_h
    port map (
            O => \N__4312\,
            I => \N__4295\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__4307\,
            I => \N__4292\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__4304\,
            I => \r_CountZ0Z_2\
        );

    \I__696\ : Odrv4
    port map (
            O => \N__4301\,
            I => \r_CountZ0Z_2\
        );

    \I__695\ : Odrv4
    port map (
            O => \N__4298\,
            I => \r_CountZ0Z_2\
        );

    \I__694\ : Odrv4
    port map (
            O => \N__4295\,
            I => \r_CountZ0Z_2\
        );

    \I__693\ : Odrv12
    port map (
            O => \N__4292\,
            I => \r_CountZ0Z_2\
        );

    \I__692\ : CascadeMux
    port map (
            O => \N__4281\,
            I => \Instance2.r_Count13_8_0_cascade_\
        );

    \I__691\ : CascadeMux
    port map (
            O => \N__4278\,
            I => \Instance2.un1_r_Count_10lt11_0_cascade_\
        );

    \I__690\ : InMux
    port map (
            O => \N__4275\,
            I => \N__4272\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__4272\,
            I => \N__4269\
        );

    \I__688\ : Odrv4
    port map (
            O => \N__4269\,
            I => \sevsegr_RNO_0Z0Z_1\
        );

    \I__687\ : InMux
    port map (
            O => \N__4266\,
            I => \N__4263\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__4263\,
            I => \r_SwitchZ0Z_3\
        );

    \I__685\ : CascadeMux
    port map (
            O => \N__4260\,
            I => \N__4257\
        );

    \I__684\ : InMux
    port map (
            O => \N__4257\,
            I => \N__4254\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__4254\,
            I => \alogicunit.m26_l_fxZ0\
        );

    \I__682\ : InMux
    port map (
            O => \N__4251\,
            I => \N__4248\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__4248\,
            I => \N__4245\
        );

    \I__680\ : Odrv4
    port map (
            O => \N__4245\,
            I => \sevsegl_RNO_0Z0Z_1\
        );

    \I__679\ : CascadeMux
    port map (
            O => \N__4242\,
            I => \N__4239\
        );

    \I__678\ : InMux
    port map (
            O => \N__4239\,
            I => \N__4235\
        );

    \I__677\ : CascadeMux
    port map (
            O => \N__4238\,
            I => \N__4232\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__4235\,
            I => \N__4227\
        );

    \I__675\ : InMux
    port map (
            O => \N__4232\,
            I => \N__4224\
        );

    \I__674\ : CascadeMux
    port map (
            O => \N__4231\,
            I => \N__4220\
        );

    \I__673\ : CascadeMux
    port map (
            O => \N__4230\,
            I => \N__4217\
        );

    \I__672\ : Span4Mux_s3_h
    port map (
            O => \N__4227\,
            I => \N__4214\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__4224\,
            I => \N__4211\
        );

    \I__670\ : InMux
    port map (
            O => \N__4223\,
            I => \N__4204\
        );

    \I__669\ : InMux
    port map (
            O => \N__4220\,
            I => \N__4204\
        );

    \I__668\ : InMux
    port map (
            O => \N__4217\,
            I => \N__4204\
        );

    \I__667\ : Odrv4
    port map (
            O => \N__4214\,
            I => \r_CountZ0Z_3\
        );

    \I__666\ : Odrv4
    port map (
            O => \N__4211\,
            I => \r_CountZ0Z_3\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__4204\,
            I => \r_CountZ0Z_3\
        );

    \I__664\ : InMux
    port map (
            O => \N__4197\,
            I => \N__4194\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__4194\,
            I => \N__4191\
        );

    \I__662\ : Odrv4
    port map (
            O => \N__4191\,
            I => \sevsegl_RNO_0Z0Z_3\
        );

    \I__661\ : InMux
    port map (
            O => \N__4188\,
            I => \N__4184\
        );

    \I__660\ : CascadeMux
    port map (
            O => \N__4187\,
            I => \N__4179\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__4184\,
            I => \N__4174\
        );

    \I__658\ : InMux
    port map (
            O => \N__4183\,
            I => \N__4171\
        );

    \I__657\ : InMux
    port map (
            O => \N__4182\,
            I => \N__4164\
        );

    \I__656\ : InMux
    port map (
            O => \N__4179\,
            I => \N__4164\
        );

    \I__655\ : InMux
    port map (
            O => \N__4178\,
            I => \N__4164\
        );

    \I__654\ : CascadeMux
    port map (
            O => \N__4177\,
            I => \N__4161\
        );

    \I__653\ : Span4Mux_s3_h
    port map (
            O => \N__4174\,
            I => \N__4157\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__4171\,
            I => \N__4154\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__4164\,
            I => \N__4151\
        );

    \I__650\ : InMux
    port map (
            O => \N__4161\,
            I => \N__4146\
        );

    \I__649\ : InMux
    port map (
            O => \N__4160\,
            I => \N__4146\
        );

    \I__648\ : Odrv4
    port map (
            O => \N__4157\,
            I => \alogicunit.result24\
        );

    \I__647\ : Odrv4
    port map (
            O => \N__4154\,
            I => \alogicunit.result24\
        );

    \I__646\ : Odrv4
    port map (
            O => \N__4151\,
            I => \alogicunit.result24\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__4146\,
            I => \alogicunit.result24\
        );

    \I__644\ : CascadeMux
    port map (
            O => \N__4137\,
            I => \alogicunit.result24_cascade_\
        );

    \I__643\ : CascadeMux
    port map (
            O => \N__4134\,
            I => \N__4130\
        );

    \I__642\ : InMux
    port map (
            O => \N__4133\,
            I => \N__4126\
        );

    \I__641\ : InMux
    port map (
            O => \N__4130\,
            I => \N__4123\
        );

    \I__640\ : InMux
    port map (
            O => \N__4129\,
            I => \N__4120\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__4126\,
            I => \N__4117\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__4123\,
            I => \N__4114\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__4120\,
            I => \alogicunit.un1_a_1_axb_3\
        );

    \I__636\ : Odrv4
    port map (
            O => \N__4117\,
            I => \alogicunit.un1_a_1_axb_3\
        );

    \I__635\ : Odrv4
    port map (
            O => \N__4114\,
            I => \alogicunit.un1_a_1_axb_3\
        );

    \I__634\ : CascadeMux
    port map (
            O => \N__4107\,
            I => \N__4103\
        );

    \I__633\ : CascadeMux
    port map (
            O => \N__4106\,
            I => \N__4100\
        );

    \I__632\ : InMux
    port map (
            O => \N__4103\,
            I => \N__4095\
        );

    \I__631\ : InMux
    port map (
            O => \N__4100\,
            I => \N__4095\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__4095\,
            I => \N__4092\
        );

    \I__629\ : Span12Mux_s3_h
    port map (
            O => \N__4092\,
            I => \N__4089\
        );

    \I__628\ : Odrv12
    port map (
            O => \N__4089\,
            I => \alogicunit.N_51\
        );

    \I__627\ : InMux
    port map (
            O => \N__4086\,
            I => \N__4080\
        );

    \I__626\ : InMux
    port map (
            O => \N__4085\,
            I => \N__4080\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__4080\,
            I => cu1_track_ns_3
        );

    \I__624\ : CascadeMux
    port map (
            O => \N__4077\,
            I => \N__4074\
        );

    \I__623\ : InMux
    port map (
            O => \N__4074\,
            I => \N__4071\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__4071\,
            I => \alogicunit.un1_a_1_cry_1_THRU_CO\
        );

    \I__621\ : InMux
    port map (
            O => \N__4068\,
            I => \alogicunit.un1_a_1_cry_1\
        );

    \I__620\ : InMux
    port map (
            O => \N__4065\,
            I => \N__4062\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__4062\,
            I => \alogicunit.un1_a_1_cry_2_THRU_CO\
        );

    \I__618\ : InMux
    port map (
            O => \N__4059\,
            I => \alogicunit.un1_a_1_cry_2\
        );

    \I__617\ : InMux
    port map (
            O => \N__4056\,
            I => \alogicunit.un1_a_1_cry_3\
        );

    \I__616\ : InMux
    port map (
            O => \N__4053\,
            I => \N__4050\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__4050\,
            I => \N__4047\
        );

    \I__614\ : Odrv4
    port map (
            O => \N__4047\,
            I => \alogicunit.result_RNO_0Z0Z_5\
        );

    \I__613\ : InMux
    port map (
            O => \N__4044\,
            I => \alogicunit.un1_a_1_cry_4\
        );

    \I__612\ : InMux
    port map (
            O => \N__4041\,
            I => \alogicunit.un1_a_1_cry_5\
        );

    \I__611\ : CascadeMux
    port map (
            O => \N__4038\,
            I => \N__4033\
        );

    \I__610\ : InMux
    port map (
            O => \N__4037\,
            I => \N__4028\
        );

    \I__609\ : InMux
    port map (
            O => \N__4036\,
            I => \N__4028\
        );

    \I__608\ : InMux
    port map (
            O => \N__4033\,
            I => \N__4025\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__4028\,
            I => \alogicunit.N_95_1\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__4025\,
            I => \alogicunit.N_95_1\
        );

    \I__605\ : InMux
    port map (
            O => \N__4020\,
            I => \alogicunit.un1_a_1_cry_6\
        );

    \I__604\ : InMux
    port map (
            O => \N__4017\,
            I => \N__4014\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__4014\,
            I => \N__4011\
        );

    \I__602\ : Odrv4
    port map (
            O => \N__4011\,
            I => left_3
        );

    \I__601\ : CascadeMux
    port map (
            O => \N__4008\,
            I => \N__4005\
        );

    \I__600\ : InMux
    port map (
            O => \N__4005\,
            I => \N__4002\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__4002\,
            I => \alogicunit.m26_l_fxZ0Z_0\
        );

    \I__598\ : CascadeMux
    port map (
            O => \N__3999\,
            I => \un1_click13_1_sn_cascade_\
        );

    \I__597\ : InMux
    port map (
            O => \N__3996\,
            I => \N__3993\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__3993\,
            I => \N__3990\
        );

    \I__595\ : Odrv12
    port map (
            O => \N__3990\,
            I => \sevsegr_RNO_0Z0Z_2\
        );

    \I__594\ : InMux
    port map (
            O => \N__3987\,
            I => \N__3984\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__3984\,
            I => \N__3979\
        );

    \I__592\ : InMux
    port map (
            O => \N__3983\,
            I => \N__3976\
        );

    \I__591\ : InMux
    port map (
            O => \N__3982\,
            I => \N__3973\
        );

    \I__590\ : Span4Mux_s3_h
    port map (
            O => \N__3979\,
            I => \N__3970\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__3976\,
            I => \r_Count11\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__3973\,
            I => \r_Count11\
        );

    \I__587\ : Odrv4
    port map (
            O => \N__3970\,
            I => \r_Count11\
        );

    \I__586\ : CascadeMux
    port map (
            O => \N__3963\,
            I => \r_Count11_cascade_\
        );

    \I__585\ : CascadeMux
    port map (
            O => \N__3960\,
            I => \alogicunit.N_95_1_cascade_\
        );

    \I__584\ : CascadeMux
    port map (
            O => \N__3957\,
            I => \N__3954\
        );

    \I__583\ : InMux
    port map (
            O => \N__3954\,
            I => \N__3951\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__3951\,
            I => \N__3948\
        );

    \I__581\ : Span4Mux_s3_h
    port map (
            O => \N__3948\,
            I => \N__3945\
        );

    \I__580\ : Odrv4
    port map (
            O => \N__3945\,
            I => right_0
        );

    \I__579\ : InMux
    port map (
            O => \N__3942\,
            I => \N__3939\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__3939\,
            I => right_3
        );

    \I__577\ : InMux
    port map (
            O => \N__3936\,
            I => \N__3933\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__3933\,
            I => \N__3930\
        );

    \I__575\ : Span4Mux_s3_h
    port map (
            O => \N__3930\,
            I => \N__3926\
        );

    \I__574\ : InMux
    port map (
            O => \N__3929\,
            I => \N__3923\
        );

    \I__573\ : Odrv4
    port map (
            O => \N__3926\,
            I => \SUM_3\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__3923\,
            I => \SUM_3\
        );

    \I__571\ : InMux
    port map (
            O => \N__3918\,
            I => \N__3915\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__3915\,
            I => \N__3912\
        );

    \I__569\ : Span4Mux_v
    port map (
            O => \N__3912\,
            I => \N__3909\
        );

    \I__568\ : Odrv4
    port map (
            O => \N__3909\,
            I => \sevsegr_RNO_1Z0Z_3\
        );

    \I__567\ : InMux
    port map (
            O => \N__3906\,
            I => \N__3903\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__3903\,
            I => \N__3900\
        );

    \I__565\ : Span4Mux_s3_h
    port map (
            O => \N__3900\,
            I => \N__3897\
        );

    \I__564\ : Odrv4
    port map (
            O => \N__3897\,
            I => right_2
        );

    \I__563\ : InMux
    port map (
            O => \N__3894\,
            I => \N__3891\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__3891\,
            I => sevsegl_7_ns_1_0
        );

    \I__561\ : InMux
    port map (
            O => \N__3888\,
            I => \N__3864\
        );

    \I__560\ : InMux
    port map (
            O => \N__3887\,
            I => \N__3864\
        );

    \I__559\ : InMux
    port map (
            O => \N__3886\,
            I => \N__3864\
        );

    \I__558\ : InMux
    port map (
            O => \N__3885\,
            I => \N__3864\
        );

    \I__557\ : InMux
    port map (
            O => \N__3884\,
            I => \N__3864\
        );

    \I__556\ : InMux
    port map (
            O => \N__3883\,
            I => \N__3864\
        );

    \I__555\ : InMux
    port map (
            O => \N__3882\,
            I => \N__3864\
        );

    \I__554\ : InMux
    port map (
            O => \N__3881\,
            I => \N__3861\
        );

    \I__553\ : InMux
    port map (
            O => \N__3880\,
            I => \N__3858\
        );

    \I__552\ : InMux
    port map (
            O => \N__3879\,
            I => \N__3855\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__3864\,
            I => \r_Switch_2_RNIK7AZ0Z11\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__3861\,
            I => \r_Switch_2_RNIK7AZ0Z11\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3858\,
            I => \r_Switch_2_RNIK7AZ0Z11\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__3855\,
            I => \r_Switch_2_RNIK7AZ0Z11\
        );

    \I__547\ : CEMux
    port map (
            O => \N__3846\,
            I => \N__3843\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__3843\,
            I => \N__3839\
        );

    \I__545\ : CEMux
    port map (
            O => \N__3842\,
            I => \N__3836\
        );

    \I__544\ : Span4Mux_h
    port map (
            O => \N__3839\,
            I => \N__3833\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__3836\,
            I => \N__3830\
        );

    \I__542\ : Odrv4
    port map (
            O => \N__3833\,
            I => un1_click17_0
        );

    \I__541\ : Odrv4
    port map (
            O => \N__3830\,
            I => un1_click17_0
        );

    \I__540\ : IoInMux
    port map (
            O => \N__3825\,
            I => \N__3822\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3822\,
            I => \r_HexEncode_i_4\
        );

    \I__538\ : IoInMux
    port map (
            O => \N__3819\,
            I => \N__3816\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__3816\,
            I => \N__3813\
        );

    \I__536\ : IoSpan4Mux
    port map (
            O => \N__3813\,
            I => \N__3810\
        );

    \I__535\ : Span4Mux_s0_v
    port map (
            O => \N__3810\,
            I => \N__3807\
        );

    \I__534\ : Odrv4
    port map (
            O => \N__3807\,
            I => \r_HexEncode_i_0\
        );

    \I__533\ : IoInMux
    port map (
            O => \N__3804\,
            I => \N__3801\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__3801\,
            I => \N__3798\
        );

    \I__531\ : IoSpan4Mux
    port map (
            O => \N__3798\,
            I => \N__3795\
        );

    \I__530\ : Odrv4
    port map (
            O => \N__3795\,
            I => \r_HexEncode_i_2\
        );

    \I__529\ : IoInMux
    port map (
            O => \N__3792\,
            I => \N__3789\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__3789\,
            I => \N__3786\
        );

    \I__527\ : IoSpan4Mux
    port map (
            O => \N__3786\,
            I => \N__3783\
        );

    \I__526\ : Odrv4
    port map (
            O => \N__3783\,
            I => \r_HexEncode_i_3\
        );

    \I__525\ : CascadeMux
    port map (
            O => \N__3780\,
            I => \N__3777\
        );

    \I__524\ : InMux
    port map (
            O => \N__3777\,
            I => \N__3774\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__3774\,
            I => \N__3765\
        );

    \I__522\ : InMux
    port map (
            O => \N__3773\,
            I => \N__3754\
        );

    \I__521\ : InMux
    port map (
            O => \N__3772\,
            I => \N__3754\
        );

    \I__520\ : InMux
    port map (
            O => \N__3771\,
            I => \N__3754\
        );

    \I__519\ : InMux
    port map (
            O => \N__3770\,
            I => \N__3754\
        );

    \I__518\ : InMux
    port map (
            O => \N__3769\,
            I => \N__3754\
        );

    \I__517\ : InMux
    port map (
            O => \N__3768\,
            I => \N__3751\
        );

    \I__516\ : Span4Mux_s1_h
    port map (
            O => \N__3765\,
            I => \N__3746\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__3754\,
            I => \N__3746\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__3751\,
            I => \sevsegrZ0Z_0\
        );

    \I__513\ : Odrv4
    port map (
            O => \N__3746\,
            I => \sevsegrZ0Z_0\
        );

    \I__512\ : InMux
    port map (
            O => \N__3741\,
            I => \N__3733\
        );

    \I__511\ : InMux
    port map (
            O => \N__3740\,
            I => \N__3722\
        );

    \I__510\ : InMux
    port map (
            O => \N__3739\,
            I => \N__3722\
        );

    \I__509\ : InMux
    port map (
            O => \N__3738\,
            I => \N__3722\
        );

    \I__508\ : InMux
    port map (
            O => \N__3737\,
            I => \N__3722\
        );

    \I__507\ : InMux
    port map (
            O => \N__3736\,
            I => \N__3722\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__3733\,
            I => \N__3716\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__3722\,
            I => \N__3716\
        );

    \I__504\ : InMux
    port map (
            O => \N__3721\,
            I => \N__3713\
        );

    \I__503\ : Odrv4
    port map (
            O => \N__3716\,
            I => \sevsegrZ0Z_2\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__3713\,
            I => \sevsegrZ0Z_2\
        );

    \I__501\ : InMux
    port map (
            O => \N__3708\,
            I => \N__3702\
        );

    \I__500\ : CascadeMux
    port map (
            O => \N__3707\,
            I => \N__3699\
        );

    \I__499\ : CascadeMux
    port map (
            O => \N__3706\,
            I => \N__3696\
        );

    \I__498\ : CascadeMux
    port map (
            O => \N__3705\,
            I => \N__3692\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3702\,
            I => \N__3688\
        );

    \I__496\ : InMux
    port map (
            O => \N__3699\,
            I => \N__3677\
        );

    \I__495\ : InMux
    port map (
            O => \N__3696\,
            I => \N__3677\
        );

    \I__494\ : InMux
    port map (
            O => \N__3695\,
            I => \N__3677\
        );

    \I__493\ : InMux
    port map (
            O => \N__3692\,
            I => \N__3677\
        );

    \I__492\ : InMux
    port map (
            O => \N__3691\,
            I => \N__3677\
        );

    \I__491\ : Sp12to4
    port map (
            O => \N__3688\,
            I => \N__3671\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__3677\,
            I => \N__3671\
        );

    \I__489\ : InMux
    port map (
            O => \N__3676\,
            I => \N__3668\
        );

    \I__488\ : Odrv12
    port map (
            O => \N__3671\,
            I => \sevsegrZ0Z_1\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__3668\,
            I => \sevsegrZ0Z_1\
        );

    \I__486\ : CascadeMux
    port map (
            O => \N__3663\,
            I => \N__3656\
        );

    \I__485\ : CascadeMux
    port map (
            O => \N__3662\,
            I => \N__3652\
        );

    \I__484\ : InMux
    port map (
            O => \N__3661\,
            I => \N__3648\
        );

    \I__483\ : InMux
    port map (
            O => \N__3660\,
            I => \N__3637\
        );

    \I__482\ : InMux
    port map (
            O => \N__3659\,
            I => \N__3637\
        );

    \I__481\ : InMux
    port map (
            O => \N__3656\,
            I => \N__3637\
        );

    \I__480\ : InMux
    port map (
            O => \N__3655\,
            I => \N__3637\
        );

    \I__479\ : InMux
    port map (
            O => \N__3652\,
            I => \N__3637\
        );

    \I__478\ : CascadeMux
    port map (
            O => \N__3651\,
            I => \N__3634\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__3648\,
            I => \N__3629\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__3637\,
            I => \N__3629\
        );

    \I__475\ : InMux
    port map (
            O => \N__3634\,
            I => \N__3626\
        );

    \I__474\ : Odrv4
    port map (
            O => \N__3629\,
            I => \sevsegrZ0Z_3\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__3626\,
            I => \sevsegrZ0Z_3\
        );

    \I__472\ : IoInMux
    port map (
            O => \N__3621\,
            I => \N__3618\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__3618\,
            I => \r_HexEncode_i_5\
        );

    \I__470\ : CascadeMux
    port map (
            O => \N__3615\,
            I => \SUM_3_cascade_\
        );

    \I__469\ : InMux
    port map (
            O => \N__3612\,
            I => \N__3609\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__3609\,
            I => \sevsegl_RNO_1Z0Z_3\
        );

    \I__467\ : InMux
    port map (
            O => \N__3606\,
            I => \N__3603\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__3603\,
            I => \N__3600\
        );

    \I__465\ : Odrv4
    port map (
            O => \N__3600\,
            I => \sevsegr_RNO_1Z0Z_1\
        );

    \I__464\ : CascadeMux
    port map (
            O => \N__3597\,
            I => \N__3594\
        );

    \I__463\ : InMux
    port map (
            O => \N__3594\,
            I => \N__3591\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__3591\,
            I => \sevsegr_RNO_1Z0Z_2\
        );

    \I__461\ : InMux
    port map (
            O => \N__3588\,
            I => \N__3585\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__3585\,
            I => \N__3582\
        );

    \I__459\ : Odrv4
    port map (
            O => \N__3582\,
            I => \sevsegr_RNO_0Z0Z_3\
        );

    \I__458\ : InMux
    port map (
            O => \N__3579\,
            I => \N__3576\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__3576\,
            I => \sevsegl_RNO_1Z0Z_1\
        );

    \I__456\ : InMux
    port map (
            O => \N__3573\,
            I => \N__3570\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__3570\,
            I => sevsegr_7_ns_1_0
        );

    \I__454\ : CascadeMux
    port map (
            O => \N__3567\,
            I => \N__3562\
        );

    \I__453\ : InMux
    port map (
            O => \N__3566\,
            I => \N__3559\
        );

    \I__452\ : InMux
    port map (
            O => \N__3565\,
            I => \N__3556\
        );

    \I__451\ : InMux
    port map (
            O => \N__3562\,
            I => \N__3553\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__3559\,
            I => \Instance1.r_CountZ0Z_14\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__3556\,
            I => \Instance1.r_CountZ0Z_14\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__3553\,
            I => \Instance1.r_CountZ0Z_14\
        );

    \I__447\ : InMux
    port map (
            O => \N__3546\,
            I => \Instance1.r_Count_2_cry_13\
        );

    \I__446\ : InMux
    port map (
            O => \N__3543\,
            I => \N__3538\
        );

    \I__445\ : InMux
    port map (
            O => \N__3542\,
            I => \N__3535\
        );

    \I__444\ : InMux
    port map (
            O => \N__3541\,
            I => \N__3532\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__3538\,
            I => \Instance1.r_CountZ0Z_15\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__3535\,
            I => \Instance1.r_CountZ0Z_15\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__3532\,
            I => \Instance1.r_CountZ0Z_15\
        );

    \I__440\ : InMux
    port map (
            O => \N__3525\,
            I => \Instance1.r_Count_2_cry_14\
        );

    \I__439\ : CascadeMux
    port map (
            O => \N__3522\,
            I => \N__3518\
        );

    \I__438\ : InMux
    port map (
            O => \N__3521\,
            I => \N__3514\
        );

    \I__437\ : InMux
    port map (
            O => \N__3518\,
            I => \N__3511\
        );

    \I__436\ : InMux
    port map (
            O => \N__3517\,
            I => \N__3508\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__3514\,
            I => \Instance1.r_CountZ0Z_16\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__3511\,
            I => \Instance1.r_CountZ0Z_16\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__3508\,
            I => \Instance1.r_CountZ0Z_16\
        );

    \I__432\ : InMux
    port map (
            O => \N__3501\,
            I => \Instance1.r_Count_2_cry_15\
        );

    \I__431\ : InMux
    port map (
            O => \N__3498\,
            I => \bfn_2_11_0_\
        );

    \I__430\ : InMux
    port map (
            O => \N__3495\,
            I => \N__3490\
        );

    \I__429\ : InMux
    port map (
            O => \N__3494\,
            I => \N__3487\
        );

    \I__428\ : InMux
    port map (
            O => \N__3493\,
            I => \N__3484\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__3490\,
            I => \Instance1.r_CountZ0Z_17\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__3487\,
            I => \Instance1.r_CountZ0Z_17\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__3484\,
            I => \Instance1.r_CountZ0Z_17\
        );

    \I__424\ : CascadeMux
    port map (
            O => \N__3477\,
            I => \N__3474\
        );

    \I__423\ : InMux
    port map (
            O => \N__3474\,
            I => \N__3468\
        );

    \I__422\ : InMux
    port map (
            O => \N__3473\,
            I => \N__3465\
        );

    \I__421\ : InMux
    port map (
            O => \N__3472\,
            I => \N__3462\
        );

    \I__420\ : InMux
    port map (
            O => \N__3471\,
            I => \N__3459\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__3468\,
            I => \N__3456\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__3465\,
            I => \Instance1.r_CountZ0Z_0\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__3462\,
            I => \Instance1.r_CountZ0Z_0\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__3459\,
            I => \Instance1.r_CountZ0Z_0\
        );

    \I__415\ : Odrv4
    port map (
            O => \N__3456\,
            I => \Instance1.r_CountZ0Z_0\
        );

    \I__414\ : SRMux
    port map (
            O => \N__3447\,
            I => \N__3435\
        );

    \I__413\ : SRMux
    port map (
            O => \N__3446\,
            I => \N__3435\
        );

    \I__412\ : SRMux
    port map (
            O => \N__3445\,
            I => \N__3435\
        );

    \I__411\ : SRMux
    port map (
            O => \N__3444\,
            I => \N__3435\
        );

    \I__410\ : GlobalMux
    port map (
            O => \N__3435\,
            I => \N__3432\
        );

    \I__409\ : gio2CtrlBuf
    port map (
            O => \N__3432\,
            I => \Instance1.r_Count12_i_g\
        );

    \I__408\ : CascadeMux
    port map (
            O => \N__3429\,
            I => \N__3426\
        );

    \I__407\ : InMux
    port map (
            O => \N__3426\,
            I => \N__3423\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__3423\,
            I => left_1
        );

    \I__405\ : CascadeMux
    port map (
            O => \N__3420\,
            I => \N__3417\
        );

    \I__404\ : InMux
    port map (
            O => \N__3417\,
            I => \N__3414\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__3414\,
            I => right_1
        );

    \I__402\ : InMux
    port map (
            O => \N__3411\,
            I => \N__3406\
        );

    \I__401\ : InMux
    port map (
            O => \N__3410\,
            I => \N__3401\
        );

    \I__400\ : InMux
    port map (
            O => \N__3409\,
            I => \N__3401\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__3406\,
            I => \Instance1.r_CountZ0Z_6\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__3401\,
            I => \Instance1.r_CountZ0Z_6\
        );

    \I__397\ : InMux
    port map (
            O => \N__3396\,
            I => \Instance1.r_Count_2_cry_5\
        );

    \I__396\ : CascadeMux
    port map (
            O => \N__3393\,
            I => \N__3388\
        );

    \I__395\ : InMux
    port map (
            O => \N__3392\,
            I => \N__3385\
        );

    \I__394\ : InMux
    port map (
            O => \N__3391\,
            I => \N__3380\
        );

    \I__393\ : InMux
    port map (
            O => \N__3388\,
            I => \N__3380\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__3385\,
            I => \N__3375\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__3380\,
            I => \N__3375\
        );

    \I__390\ : Odrv4
    port map (
            O => \N__3375\,
            I => \Instance1.r_CountZ0Z_7\
        );

    \I__389\ : InMux
    port map (
            O => \N__3372\,
            I => \Instance1.r_Count_2_cry_6\
        );

    \I__388\ : InMux
    port map (
            O => \N__3369\,
            I => \N__3364\
        );

    \I__387\ : InMux
    port map (
            O => \N__3368\,
            I => \N__3359\
        );

    \I__386\ : InMux
    port map (
            O => \N__3367\,
            I => \N__3359\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__3364\,
            I => \Instance1.r_CountZ0Z_8\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__3359\,
            I => \Instance1.r_CountZ0Z_8\
        );

    \I__383\ : InMux
    port map (
            O => \N__3354\,
            I => \Instance1.r_Count_2_cry_7\
        );

    \I__382\ : CascadeMux
    port map (
            O => \N__3351\,
            I => \N__3346\
        );

    \I__381\ : InMux
    port map (
            O => \N__3350\,
            I => \N__3343\
        );

    \I__380\ : InMux
    port map (
            O => \N__3349\,
            I => \N__3340\
        );

    \I__379\ : InMux
    port map (
            O => \N__3346\,
            I => \N__3337\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__3343\,
            I => \Instance1.r_CountZ0Z_9\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__3340\,
            I => \Instance1.r_CountZ0Z_9\
        );

    \I__376\ : LocalMux
    port map (
            O => \N__3337\,
            I => \Instance1.r_CountZ0Z_9\
        );

    \I__375\ : InMux
    port map (
            O => \N__3330\,
            I => \bfn_2_10_0_\
        );

    \I__374\ : CascadeMux
    port map (
            O => \N__3327\,
            I => \N__3324\
        );

    \I__373\ : InMux
    port map (
            O => \N__3324\,
            I => \N__3319\
        );

    \I__372\ : InMux
    port map (
            O => \N__3323\,
            I => \N__3316\
        );

    \I__371\ : InMux
    port map (
            O => \N__3322\,
            I => \N__3313\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__3319\,
            I => \Instance1.r_CountZ0Z_10\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__3316\,
            I => \Instance1.r_CountZ0Z_10\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__3313\,
            I => \Instance1.r_CountZ0Z_10\
        );

    \I__367\ : InMux
    port map (
            O => \N__3306\,
            I => \Instance1.r_Count_2_cry_9\
        );

    \I__366\ : InMux
    port map (
            O => \N__3303\,
            I => \N__3298\
        );

    \I__365\ : InMux
    port map (
            O => \N__3302\,
            I => \N__3295\
        );

    \I__364\ : InMux
    port map (
            O => \N__3301\,
            I => \N__3292\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__3298\,
            I => \Instance1.r_CountZ0Z_11\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__3295\,
            I => \Instance1.r_CountZ0Z_11\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__3292\,
            I => \Instance1.r_CountZ0Z_11\
        );

    \I__360\ : InMux
    port map (
            O => \N__3285\,
            I => \Instance1.r_Count_2_cry_10\
        );

    \I__359\ : CascadeMux
    port map (
            O => \N__3282\,
            I => \N__3278\
        );

    \I__358\ : InMux
    port map (
            O => \N__3281\,
            I => \N__3274\
        );

    \I__357\ : InMux
    port map (
            O => \N__3278\,
            I => \N__3269\
        );

    \I__356\ : InMux
    port map (
            O => \N__3277\,
            I => \N__3269\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__3274\,
            I => \Instance1.r_CountZ0Z_12\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__3269\,
            I => \Instance1.r_CountZ0Z_12\
        );

    \I__353\ : InMux
    port map (
            O => \N__3264\,
            I => \Instance1.r_Count_2_cry_11\
        );

    \I__352\ : InMux
    port map (
            O => \N__3261\,
            I => \N__3256\
        );

    \I__351\ : InMux
    port map (
            O => \N__3260\,
            I => \N__3251\
        );

    \I__350\ : InMux
    port map (
            O => \N__3259\,
            I => \N__3251\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__3256\,
            I => \Instance1.r_CountZ0Z_13\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__3251\,
            I => \Instance1.r_CountZ0Z_13\
        );

    \I__347\ : InMux
    port map (
            O => \N__3246\,
            I => \Instance1.r_Count_2_cry_12\
        );

    \I__346\ : CascadeMux
    port map (
            O => \N__3243\,
            I => \SUM_2_cascade_\
        );

    \I__345\ : IoInMux
    port map (
            O => \N__3240\,
            I => \N__3237\
        );

    \I__344\ : LocalMux
    port map (
            O => \N__3237\,
            I => \r_HexEncode_i_0_0\
        );

    \I__343\ : IoInMux
    port map (
            O => \N__3234\,
            I => \N__3231\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__3231\,
            I => \r_HexEncode_i_0_1\
        );

    \I__341\ : IoInMux
    port map (
            O => \N__3228\,
            I => \N__3225\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__3225\,
            I => \r_HexEncode_i_6\
        );

    \I__339\ : InMux
    port map (
            O => \N__3222\,
            I => \N__3217\
        );

    \I__338\ : InMux
    port map (
            O => \N__3221\,
            I => \N__3212\
        );

    \I__337\ : InMux
    port map (
            O => \N__3220\,
            I => \N__3212\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__3217\,
            I => \Instance1.r_CountZ0Z_1\
        );

    \I__335\ : LocalMux
    port map (
            O => \N__3212\,
            I => \Instance1.r_CountZ0Z_1\
        );

    \I__334\ : InMux
    port map (
            O => \N__3207\,
            I => \N__3203\
        );

    \I__333\ : InMux
    port map (
            O => \N__3206\,
            I => \N__3200\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__3203\,
            I => \Instance1.r_CountZ0Z_2\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__3200\,
            I => \Instance1.r_CountZ0Z_2\
        );

    \I__330\ : InMux
    port map (
            O => \N__3195\,
            I => \Instance1.r_Count_2_cry_1\
        );

    \I__329\ : CascadeMux
    port map (
            O => \N__3192\,
            I => \N__3188\
        );

    \I__328\ : InMux
    port map (
            O => \N__3191\,
            I => \N__3185\
        );

    \I__327\ : InMux
    port map (
            O => \N__3188\,
            I => \N__3182\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__3185\,
            I => \Instance1.r_CountZ0Z_3\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__3182\,
            I => \Instance1.r_CountZ0Z_3\
        );

    \I__324\ : InMux
    port map (
            O => \N__3177\,
            I => \Instance1.r_Count_2_cry_2\
        );

    \I__323\ : InMux
    port map (
            O => \N__3174\,
            I => \N__3169\
        );

    \I__322\ : InMux
    port map (
            O => \N__3173\,
            I => \N__3166\
        );

    \I__321\ : InMux
    port map (
            O => \N__3172\,
            I => \N__3163\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__3169\,
            I => \N__3158\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__3166\,
            I => \N__3158\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__3163\,
            I => \Instance1.r_CountZ0Z_4\
        );

    \I__317\ : Odrv12
    port map (
            O => \N__3158\,
            I => \Instance1.r_CountZ0Z_4\
        );

    \I__316\ : InMux
    port map (
            O => \N__3153\,
            I => \Instance1.r_Count_2_cry_3\
        );

    \I__315\ : InMux
    port map (
            O => \N__3150\,
            I => \N__3147\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__3147\,
            I => \N__3142\
        );

    \I__313\ : InMux
    port map (
            O => \N__3146\,
            I => \N__3139\
        );

    \I__312\ : InMux
    port map (
            O => \N__3145\,
            I => \N__3136\
        );

    \I__311\ : Odrv4
    port map (
            O => \N__3142\,
            I => \Instance1.r_CountZ0Z_5\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__3139\,
            I => \Instance1.r_CountZ0Z_5\
        );

    \I__309\ : LocalMux
    port map (
            O => \N__3136\,
            I => \Instance1.r_CountZ0Z_5\
        );

    \I__308\ : InMux
    port map (
            O => \N__3129\,
            I => \Instance1.r_Count_2_cry_4\
        );

    \I__307\ : CascadeMux
    port map (
            O => \N__3126\,
            I => \sevsegl_RNO_0Z0Z_2_cascade_\
        );

    \I__306\ : InMux
    port map (
            O => \N__3123\,
            I => \N__3120\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__3120\,
            I => \sevsegl_RNO_1Z0Z_2\
        );

    \I__304\ : IoInMux
    port map (
            O => \N__3117\,
            I => \N__3114\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__3114\,
            I => \r_HexEncode_i_0_6\
        );

    \I__302\ : IoInMux
    port map (
            O => \N__3111\,
            I => \N__3108\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__3108\,
            I => \r_HexEncode_i_1\
        );

    \I__300\ : IoInMux
    port map (
            O => \N__3105\,
            I => \N__3102\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__3102\,
            I => \r_HexEncode_i_0_5\
        );

    \I__298\ : InMux
    port map (
            O => \N__3099\,
            I => \N__3096\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__3096\,
            I => \SUM_2\
        );

    \I__296\ : InMux
    port map (
            O => \N__3093\,
            I => \N__3090\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__3090\,
            I => \Instance1.un1_r_Count_10lto17_1\
        );

    \I__294\ : InMux
    port map (
            O => \N__3087\,
            I => \N__3084\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__3084\,
            I => \r_SwitchZ0Z_1\
        );

    \I__292\ : InMux
    port map (
            O => \N__3081\,
            I => \N__3078\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__3078\,
            I => \N__3075\
        );

    \I__290\ : Odrv4
    port map (
            O => \N__3075\,
            I => \Instance1.r_Count13_8_0\
        );

    \I__289\ : CascadeMux
    port map (
            O => \N__3072\,
            I => \Instance1.r_Count13_4_cascade_\
        );

    \I__288\ : InMux
    port map (
            O => \N__3069\,
            I => \N__3066\
        );

    \I__287\ : LocalMux
    port map (
            O => \N__3066\,
            I => \Instance1.r_Count13_7\
        );

    \I__286\ : InMux
    port map (
            O => \N__3063\,
            I => \N__3060\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__3060\,
            I => \N__3057\
        );

    \I__284\ : Odrv4
    port map (
            O => \N__3057\,
            I => \Instance1.r_Count13_10\
        );

    \I__283\ : InMux
    port map (
            O => \N__3054\,
            I => \N__3050\
        );

    \I__282\ : InMux
    port map (
            O => \N__3053\,
            I => \N__3047\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__3050\,
            I => \N__3044\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__3047\,
            I => \N__3041\
        );

    \I__279\ : Span4Mux_v
    port map (
            O => \N__3044\,
            I => \N__3038\
        );

    \I__278\ : Sp12to4
    port map (
            O => \N__3041\,
            I => \N__3033\
        );

    \I__277\ : Sp12to4
    port map (
            O => \N__3038\,
            I => \N__3033\
        );

    \I__276\ : Span12Mux_v
    port map (
            O => \N__3033\,
            I => \N__3030\
        );

    \I__275\ : Odrv12
    port map (
            O => \N__3030\,
            I => \i_Switch_1_c\
        );

    \I__274\ : InMux
    port map (
            O => \N__3027\,
            I => \N__3024\
        );

    \I__273\ : LocalMux
    port map (
            O => \N__3024\,
            I => \Instance1.r_Count13_12\
        );

    \I__272\ : CascadeMux
    port map (
            O => \N__3021\,
            I => \Instance1.r_Count13_13_cascade_\
        );

    \I__271\ : InMux
    port map (
            O => \N__3018\,
            I => \N__3015\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__3015\,
            I => \N__3009\
        );

    \I__269\ : InMux
    port map (
            O => \N__3014\,
            I => \N__3002\
        );

    \I__268\ : InMux
    port map (
            O => \N__3013\,
            I => \N__3002\
        );

    \I__267\ : InMux
    port map (
            O => \N__3012\,
            I => \N__3002\
        );

    \I__266\ : Odrv12
    port map (
            O => \N__3009\,
            I => \w_Switch_1\
        );

    \I__265\ : LocalMux
    port map (
            O => \N__3002\,
            I => \w_Switch_1\
        );

    \I__264\ : CascadeMux
    port map (
            O => \N__2997\,
            I => \Instance1.un1_r_Count_10lt11_0_cascade_\
        );

    \I__263\ : InMux
    port map (
            O => \N__2994\,
            I => \N__2991\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__2991\,
            I => \Instance1.un1_r_Count_10lto11_1\
        );

    \I__261\ : CascadeMux
    port map (
            O => \N__2988\,
            I => \Instance1.un1_r_Count_10lt17_cascade_\
        );

    \I__260\ : IoInMux
    port map (
            O => \N__2985\,
            I => \N__2982\
        );

    \I__259\ : LocalMux
    port map (
            O => \N__2982\,
            I => \Instance1.r_Count12_i\
        );

    \IN_MUX_bfv_4_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_12_0_\
        );

    \IN_MUX_bfv_6_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_7_0_\
        );

    \IN_MUX_bfv_6_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Instance4.r_Count_2_cry_8\,
            carryinitout => \bfn_6_8_0_\
        );

    \IN_MUX_bfv_6_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Instance4.r_Count_2_cry_16\,
            carryinitout => \bfn_6_9_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Instance3.r_Count_2_cry_8\,
            carryinitout => \bfn_8_10_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Instance3.r_Count_2_cry_16\,
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_6_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_10_0_\
        );

    \IN_MUX_bfv_6_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Instance2.r_Count_2_cry_8\,
            carryinitout => \bfn_6_11_0_\
        );

    \IN_MUX_bfv_6_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Instance2.r_Count_2_cry_16\,
            carryinitout => \bfn_6_12_0_\
        );

    \IN_MUX_bfv_2_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_9_0_\
        );

    \IN_MUX_bfv_2_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Instance1.r_Count_2_cry_8\,
            carryinitout => \bfn_2_10_0_\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Instance1.r_Count_2_cry_16\,
            carryinitout => \bfn_2_11_0_\
        );

    \Instance1.r_State_RNIK9757_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2985\,
            GLOBALBUFFEROUTPUT => \Instance1.r_Count12_i_g\
        );

    \Instance4.r_State_RNI4ONP3_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__6204\,
            GLOBALBUFFEROUTPUT => \Instance4.r_Count12_i_g\
        );

    \Instance2.r_State_RNI4PC15_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4839\,
            GLOBALBUFFEROUTPUT => \Instance2.r_Count12_i_g\
        );

    \Instance3.r_State_RNIK8IT5_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__6498\,
            GLOBALBUFFEROUTPUT => \Instance3.r_Count12_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \Instance1.r_State_RNO_5_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__3410\,
            in1 => \N__3542\,
            in2 => \N__3522\,
            in3 => \N__3368\,
            lcout => \Instance1.r_Count13_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance1.r_Count_RNIC2TU1_8_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3322\,
            in1 => \N__3301\,
            in2 => \N__3351\,
            in3 => \N__3367\,
            lcout => \Instance1.un1_r_Count_10lto11_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance1.r_Count_RNIED2U1_4_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__3173\,
            in1 => \N__3145\,
            in2 => \N__3393\,
            in3 => \N__3409\,
            lcout => OPEN,
            ltout => \Instance1.un1_r_Count_10lt11_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance1.r_Count_RNID9RS4_12_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100010001"
        )
    port map (
            in0 => \N__3277\,
            in1 => \N__3259\,
            in2 => \N__2997\,
            in3 => \N__2994\,
            lcout => OPEN,
            ltout => \Instance1.un1_r_Count_10lt17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance1.r_State_RNIK9757_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111110011001"
        )
    port map (
            in0 => \N__3054\,
            in1 => \N__3018\,
            in2 => \N__2988\,
            in3 => \N__3093\,
            lcout => \Instance1.r_Count12_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance1.r_State_RNO_3_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__3174\,
            in1 => \N__3391\,
            in2 => \N__3282\,
            in3 => \N__3260\,
            lcout => \Instance1.r_Count13_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance1.r_Count_RNIIVNV1_17_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3493\,
            in1 => \N__3541\,
            in2 => \N__3567\,
            in3 => \N__3517\,
            lcout => \Instance1.un1_r_Count_10lto17_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance1.r_State_RNO_4_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3206\,
            in1 => \N__3220\,
            in2 => \N__3192\,
            in3 => \N__3350\,
            lcout => \Instance1.r_Count13_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance1.r_Count_1_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__3221\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3473\,
            lcout => \Instance1.r_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7081\,
            ce => 'H',
            sr => \N__3444\
        );

    \r_Switch_1_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__3014\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \r_SwitchZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7083\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance1.r_State_RNIPV6C_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3087\,
            in2 => \_gnd_net_\,
            in3 => \N__3012\,
            lcout => click13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance1.r_State_RNO_2_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3565\,
            in2 => \_gnd_net_\,
            in3 => \N__3494\,
            lcout => OPEN,
            ltout => \Instance1.r_Count13_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance1.r_State_RNO_0_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__3471\,
            in1 => \N__3081\,
            in2 => \N__3072\,
            in3 => \N__3150\,
            lcout => \Instance1.r_Count13_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance1.r_State_RNO_1_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__3069\,
            in1 => \N__3303\,
            in2 => \N__3327\,
            in3 => \N__3063\,
            lcout => OPEN,
            ltout => \Instance1.r_Count13_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance1.r_State_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__3053\,
            in1 => \N__3027\,
            in2 => \N__3021\,
            in3 => \N__3013\,
            lcout => \w_Switch_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7083\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance2.r_State_RNIHFHJ2_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__4579\,
            in1 => \N__3987\,
            in2 => \_gnd_net_\,
            in3 => \N__4761\,
            lcout => un1_click17_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_Switch_2_RNIK7A11_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__4917\,
            in1 => \N__4578\,
            in2 => \_gnd_net_\,
            in3 => \N__4833\,
            lcout => \r_Switch_2_RNIK7AZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sevsegl_RNO_0_2_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__4332\,
            in1 => \N__4527\,
            in2 => \_gnd_net_\,
            in3 => \N__4806\,
            lcout => OPEN,
            ltout => \sevsegl_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sevsegl_2_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3123\,
            in2 => \N__3126\,
            in3 => \N__3881\,
            lcout => \sevseglZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7085\,
            ce => \N__3842\,
            sr => \_gnd_net_\
        );

    \sevsegl_RNO_1_2_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4710\,
            in1 => \N__3099\,
            in2 => \_gnd_net_\,
            in3 => \N__4604\,
            lcout => \sevsegl_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sevsegr_RNO_0_0_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100101110"
        )
    port map (
            in0 => \N__4386\,
            in1 => \N__4809\,
            in2 => \N__4491\,
            in3 => \N__3880\,
            lcout => sevsegr_7_ns_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SegInst1.r_HexEncode_i_6_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000100000010"
        )
    port map (
            in0 => \N__6060\,
            in1 => \N__6017\,
            in2 => \N__5970\,
            in3 => \N__5913\,
            lcout => \r_HexEncode_i_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7088\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SegInst2.r_HexEncode_i_1_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010110100000100"
        )
    port map (
            in0 => \N__3721\,
            in1 => \N__3676\,
            in2 => \N__3651\,
            in3 => \N__3768\,
            lcout => \r_HexEncode_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7088\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SegInst1.r_HexEncode_i_5_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001010101000"
        )
    port map (
            in0 => \N__6059\,
            in1 => \N__6016\,
            in2 => \N__5969\,
            in3 => \N__5912\,
            lcout => \r_HexEncode_i_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7088\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance2.SUM_2_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__4331\,
            in1 => \N__4454\,
            in2 => \_gnd_net_\,
            in3 => \N__4385\,
            lcout => \SUM_2\,
            ltout => \SUM_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sevsegr_RNO_1_2_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__4605\,
            in1 => \_gnd_net_\,
            in2 => \N__3243\,
            in3 => \N__3906\,
            lcout => \sevsegr_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SegInst1.r_HexEncode_iZ0Z_0_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100100100001"
        )
    port map (
            in0 => \N__6066\,
            in1 => \N__6018\,
            in2 => \N__5971\,
            in3 => \N__5914\,
            lcout => \r_HexEncode_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7092\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SegInst1.r_HexEncode_i_1_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100000110010"
        )
    port map (
            in0 => \N__5915\,
            in1 => \N__5963\,
            in2 => \N__6030\,
            in3 => \N__6067\,
            lcout => \r_HexEncode_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7092\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SegInst2.r_HexEncode_i_6_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000000010100"
        )
    port map (
            in0 => \N__3708\,
            in1 => \N__3741\,
            in2 => \N__3780\,
            in3 => \N__3661\,
            lcout => \r_HexEncode_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7102\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance1.r_Count_2_cry_1_c_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3222\,
            in2 => \N__3477\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_9_0_\,
            carryout => \Instance1.r_Count_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance1.r_Count_2_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3207\,
            in2 => \_gnd_net_\,
            in3 => \N__3195\,
            lcout => \Instance1.r_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \Instance1.r_Count_2_cry_1\,
            carryout => \Instance1.r_Count_2_cry_2\,
            clk => \N__7082\,
            ce => 'H',
            sr => \N__3445\
        );

    \Instance1.r_Count_3_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3191\,
            in2 => \_gnd_net_\,
            in3 => \N__3177\,
            lcout => \Instance1.r_CountZ0Z_3\,
            ltout => OPEN,
            carryin => \Instance1.r_Count_2_cry_2\,
            carryout => \Instance1.r_Count_2_cry_3\,
            clk => \N__7082\,
            ce => 'H',
            sr => \N__3445\
        );

    \Instance1.r_Count_4_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3172\,
            in2 => \_gnd_net_\,
            in3 => \N__3153\,
            lcout => \Instance1.r_CountZ0Z_4\,
            ltout => OPEN,
            carryin => \Instance1.r_Count_2_cry_3\,
            carryout => \Instance1.r_Count_2_cry_4\,
            clk => \N__7082\,
            ce => 'H',
            sr => \N__3445\
        );

    \Instance1.r_Count_5_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3146\,
            in2 => \_gnd_net_\,
            in3 => \N__3129\,
            lcout => \Instance1.r_CountZ0Z_5\,
            ltout => OPEN,
            carryin => \Instance1.r_Count_2_cry_4\,
            carryout => \Instance1.r_Count_2_cry_5\,
            clk => \N__7082\,
            ce => 'H',
            sr => \N__3445\
        );

    \Instance1.r_Count_6_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3411\,
            in2 => \_gnd_net_\,
            in3 => \N__3396\,
            lcout => \Instance1.r_CountZ0Z_6\,
            ltout => OPEN,
            carryin => \Instance1.r_Count_2_cry_5\,
            carryout => \Instance1.r_Count_2_cry_6\,
            clk => \N__7082\,
            ce => 'H',
            sr => \N__3445\
        );

    \Instance1.r_Count_7_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3392\,
            in2 => \_gnd_net_\,
            in3 => \N__3372\,
            lcout => \Instance1.r_CountZ0Z_7\,
            ltout => OPEN,
            carryin => \Instance1.r_Count_2_cry_6\,
            carryout => \Instance1.r_Count_2_cry_7\,
            clk => \N__7082\,
            ce => 'H',
            sr => \N__3445\
        );

    \Instance1.r_Count_8_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3369\,
            in2 => \_gnd_net_\,
            in3 => \N__3354\,
            lcout => \Instance1.r_CountZ0Z_8\,
            ltout => OPEN,
            carryin => \Instance1.r_Count_2_cry_7\,
            carryout => \Instance1.r_Count_2_cry_8\,
            clk => \N__7082\,
            ce => 'H',
            sr => \N__3445\
        );

    \Instance1.r_Count_9_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3349\,
            in2 => \_gnd_net_\,
            in3 => \N__3330\,
            lcout => \Instance1.r_CountZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_2_10_0_\,
            carryout => \Instance1.r_Count_2_cry_9\,
            clk => \N__7084\,
            ce => 'H',
            sr => \N__3446\
        );

    \Instance1.r_Count_10_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3323\,
            in2 => \_gnd_net_\,
            in3 => \N__3306\,
            lcout => \Instance1.r_CountZ0Z_10\,
            ltout => OPEN,
            carryin => \Instance1.r_Count_2_cry_9\,
            carryout => \Instance1.r_Count_2_cry_10\,
            clk => \N__7084\,
            ce => 'H',
            sr => \N__3446\
        );

    \Instance1.r_Count_11_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3302\,
            in2 => \_gnd_net_\,
            in3 => \N__3285\,
            lcout => \Instance1.r_CountZ0Z_11\,
            ltout => OPEN,
            carryin => \Instance1.r_Count_2_cry_10\,
            carryout => \Instance1.r_Count_2_cry_11\,
            clk => \N__7084\,
            ce => 'H',
            sr => \N__3446\
        );

    \Instance1.r_Count_12_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3281\,
            in2 => \_gnd_net_\,
            in3 => \N__3264\,
            lcout => \Instance1.r_CountZ0Z_12\,
            ltout => OPEN,
            carryin => \Instance1.r_Count_2_cry_11\,
            carryout => \Instance1.r_Count_2_cry_12\,
            clk => \N__7084\,
            ce => 'H',
            sr => \N__3446\
        );

    \Instance1.r_Count_13_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3261\,
            in2 => \_gnd_net_\,
            in3 => \N__3246\,
            lcout => \Instance1.r_CountZ0Z_13\,
            ltout => OPEN,
            carryin => \Instance1.r_Count_2_cry_12\,
            carryout => \Instance1.r_Count_2_cry_13\,
            clk => \N__7084\,
            ce => 'H',
            sr => \N__3446\
        );

    \Instance1.r_Count_14_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3566\,
            in2 => \_gnd_net_\,
            in3 => \N__3546\,
            lcout => \Instance1.r_CountZ0Z_14\,
            ltout => OPEN,
            carryin => \Instance1.r_Count_2_cry_13\,
            carryout => \Instance1.r_Count_2_cry_14\,
            clk => \N__7084\,
            ce => 'H',
            sr => \N__3446\
        );

    \Instance1.r_Count_15_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3543\,
            in2 => \_gnd_net_\,
            in3 => \N__3525\,
            lcout => \Instance1.r_CountZ0Z_15\,
            ltout => OPEN,
            carryin => \Instance1.r_Count_2_cry_14\,
            carryout => \Instance1.r_Count_2_cry_15\,
            clk => \N__7084\,
            ce => 'H',
            sr => \N__3446\
        );

    \Instance1.r_Count_16_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3521\,
            in2 => \_gnd_net_\,
            in3 => \N__3501\,
            lcout => \Instance1.r_CountZ0Z_16\,
            ltout => OPEN,
            carryin => \Instance1.r_Count_2_cry_15\,
            carryout => \Instance1.r_Count_2_cry_16\,
            clk => \N__7084\,
            ce => 'H',
            sr => \N__3446\
        );

    \Instance1.r_Count_17_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3495\,
            in2 => \_gnd_net_\,
            in3 => \N__3498\,
            lcout => \Instance1.r_CountZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7086\,
            ce => 'H',
            sr => \N__3447\
        );

    \Instance1.r_Count_0_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3472\,
            lcout => \Instance1.r_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7086\,
            ce => 'H',
            sr => \N__3447\
        );

    \alogicunit.result_1_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__4508\,
            in1 => \N__4188\,
            in2 => \N__4106\,
            in3 => \N__5147\,
            lcout => right_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7089\,
            ce => \N__5405\,
            sr => \_gnd_net_\
        );

    \alogicunit.result_5_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__4509\,
            in1 => \N__5148\,
            in2 => \N__4107\,
            in3 => \N__4053\,
            lcout => left_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7089\,
            ce => \N__5405\,
            sr => \_gnd_net_\
        );

    \sevsegl_RNO_1_1_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__4388\,
            in1 => \N__4460\,
            in2 => \N__3429\,
            in3 => \N__4580\,
            lcout => \sevsegl_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sevsegr_RNO_1_1_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__4581\,
            in1 => \N__4459\,
            in2 => \N__3420\,
            in3 => \N__4387\,
            lcout => \sevsegr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sevsegl_RNO_1_3_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4017\,
            in1 => \N__3936\,
            in2 => \_gnd_net_\,
            in3 => \N__4582\,
            lcout => \sevsegl_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sevsegr_RNO_0_3_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__4807\,
            in1 => \N__5337\,
            in2 => \N__4242\,
            in3 => \N__5146\,
            lcout => \sevsegr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sevsegl_RNO_0_0_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100101110"
        )
    port map (
            in0 => \N__4389\,
            in1 => \N__4808\,
            in2 => \N__4490\,
            in3 => \N__3879\,
            lcout => sevsegl_7_ns_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sevsegl_3_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__3884\,
            in1 => \N__4197\,
            in2 => \_gnd_net_\,
            in3 => \N__3612\,
            lcout => \sevseglZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7093\,
            ce => \N__3846\,
            sr => \_gnd_net_\
        );

    \sevsegr_1_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__3606\,
            in1 => \N__4275\,
            in2 => \_gnd_net_\,
            in3 => \N__3886\,
            lcout => \sevsegrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7093\,
            ce => \N__3846\,
            sr => \_gnd_net_\
        );

    \sevsegr_2_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__3887\,
            in1 => \_gnd_net_\,
            in2 => \N__3597\,
            in3 => \N__3996\,
            lcout => \sevsegrZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7093\,
            ce => \N__3846\,
            sr => \_gnd_net_\
        );

    \sevsegr_3_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3588\,
            in1 => \N__3918\,
            in2 => \_gnd_net_\,
            in3 => \N__3888\,
            lcout => \sevsegrZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7093\,
            ce => \N__3846\,
            sr => \_gnd_net_\
        );

    \sevsegl_1_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__3883\,
            in1 => \N__3579\,
            in2 => \_gnd_net_\,
            in3 => \N__4251\,
            lcout => \sevseglZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7093\,
            ce => \N__3846\,
            sr => \_gnd_net_\
        );

    \sevsegr_0_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__3573\,
            in1 => \N__4621\,
            in2 => \N__3957\,
            in3 => \N__3885\,
            lcout => \sevsegrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7093\,
            ce => \N__3846\,
            sr => \_gnd_net_\
        );

    \sevsegl_0_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__3894\,
            in1 => \N__4620\,
            in2 => \N__4740\,
            in3 => \N__3882\,
            lcout => \sevseglZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7093\,
            ce => \N__3846\,
            sr => \_gnd_net_\
        );

    \SegInst2.r_HexEncode_i_4_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010000010000"
        )
    port map (
            in0 => \N__3770\,
            in1 => \N__3739\,
            in2 => \N__3706\,
            in3 => \N__3659\,
            lcout => \r_HexEncode_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SegInst2.r_HexEncode_i_0_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100100100001"
        )
    port map (
            in0 => \N__3736\,
            in1 => \N__3691\,
            in2 => \N__3662\,
            in3 => \N__3772\,
            lcout => \r_HexEncode_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SegInst2.r_HexEncode_i_2_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001010101110"
        )
    port map (
            in0 => \N__3769\,
            in1 => \N__3737\,
            in2 => \N__3705\,
            in3 => \N__3655\,
            lcout => \r_HexEncode_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SegInst2.r_HexEncode_i_3_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100101000010"
        )
    port map (
            in0 => \N__3738\,
            in1 => \N__3695\,
            in2 => \N__3663\,
            in3 => \N__3773\,
            lcout => \r_HexEncode_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SegInst2.r_HexEncode_i_5_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001001000"
        )
    port map (
            in0 => \N__3771\,
            in1 => \N__3740\,
            in2 => \N__3707\,
            in3 => \N__3660\,
            lcout => \r_HexEncode_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_Count_1_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001011110000"
        )
    port map (
            in0 => \N__4362\,
            in1 => \N__3982\,
            in2 => \N__4438\,
            in3 => \N__4623\,
            lcout => \r_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7090\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance2.SUM_3_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__4322\,
            in1 => \N__4419\,
            in2 => \N__4230\,
            in3 => \N__4359\,
            lcout => \SUM_3\,
            ltout => \SUM_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_Count_3_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__3983\,
            in1 => \N__4223\,
            in2 => \N__3615\,
            in3 => \N__4624\,
            lcout => \r_CountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7090\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance2.r_Count11_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__4323\,
            in1 => \N__4418\,
            in2 => \N__4231\,
            in3 => \N__4360\,
            lcout => \r_Count11\,
            ltout => \r_Count11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_Count_0_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010110101010"
        )
    port map (
            in0 => \N__4361\,
            in1 => \_gnd_net_\,
            in2 => \N__3963\,
            in3 => \N__4622\,
            lcout => \r_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7090\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alogicunit.result_13_iv_3_140_i_a4_1_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000101"
        )
    port map (
            in0 => \N__5143\,
            in1 => \N__5327\,
            in2 => \N__5234\,
            in3 => \N__5038\,
            lcout => \alogicunit.N_95_1\,
            ltout => \alogicunit.N_95_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alogicunit.result_0_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3960\,
            in3 => \N__4643\,
            lcout => right_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7094\,
            ce => \N__5406\,
            sr => \_gnd_net_\
        );

    \alogicunit.result_3_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010011111000"
        )
    port map (
            in0 => \N__4133\,
            in1 => \N__4037\,
            in2 => \N__4647\,
            in3 => \N__4065\,
            lcout => right_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7094\,
            ce => \N__5406\,
            sr => \_gnd_net_\
        );

    \sevsegr_RNO_1_3_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__4606\,
            in1 => \N__3942\,
            in2 => \_gnd_net_\,
            in3 => \N__3929\,
            lcout => \sevsegr_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alogicunit.result_2_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111011101010"
        )
    port map (
            in0 => \N__4539\,
            in1 => \N__4036\,
            in2 => \N__4077\,
            in3 => \N__4183\,
            lcout => right_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7094\,
            ce => \N__5406\,
            sr => \_gnd_net_\
        );

    \alogicunit.negative_e_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__5144\,
            in1 => \N__5328\,
            in2 => \N__5235\,
            in3 => \N__5039\,
            lcout => negative,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7094\,
            ce => \N__5406\,
            sr => \_gnd_net_\
        );

    \alogicunit.un1_a_1_cry_1_c_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4697\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_12_0_\,
            carryout => \alogicunit.un1_a_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alogicunit.un1_a_1_cry_1_THRU_LUT4_0_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4178\,
            in2 => \_gnd_net_\,
            in3 => \N__4068\,
            lcout => \alogicunit.un1_a_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \alogicunit.un1_a_1_cry_1\,
            carryout => \alogicunit.un1_a_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alogicunit.un1_a_1_cry_2_THRU_LUT4_0_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4134\,
            in3 => \N__4059\,
            lcout => \alogicunit.un1_a_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \alogicunit.un1_a_1_cry_2\,
            carryout => \alogicunit.un1_a_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alogicunit.result_RNO_0_4_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5363\,
            in2 => \N__4008\,
            in3 => \N__4056\,
            lcout => \alogicunit.result_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \alogicunit.un1_a_1_cry_3\,
            carryout => \alogicunit.un1_a_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alogicunit.result_RNO_0_5_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6105\,
            in2 => \N__4187\,
            in3 => \N__4044\,
            lcout => \alogicunit.result_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \alogicunit.un1_a_1_cry_4\,
            carryout => \alogicunit.un1_a_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alogicunit.result_RNO_0_6_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5364\,
            in2 => \N__4260\,
            in3 => \N__4041\,
            lcout => \alogicunit.result_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \alogicunit.un1_a_1_cry_5\,
            carryout => \alogicunit.un1_a_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alogicunit.result_7_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110011101100"
        )
    port map (
            in0 => \N__4182\,
            in1 => \N__4538\,
            in2 => \N__4038\,
            in3 => \N__4020\,
            lcout => left_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7098\,
            ce => \N__5404\,
            sr => \_gnd_net_\
        );

    \alogicunit.m26_l_fx_0_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5356\,
            in2 => \_gnd_net_\,
            in3 => \N__4160\,
            lcout => \alogicunit.m26_l_fxZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance2.un1_w_Switch_3_1_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6555\,
            in2 => \_gnd_net_\,
            in3 => \N__4266\,
            lcout => un1_click13_1_sn,
            ltout => \un1_click13_1_sn_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sevsegr_RNO_0_2_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4327\,
            in2 => \N__3999\,
            in3 => \N__4520\,
            lcout => \sevsegr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sevsegr_RNO_0_1_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010101100"
        )
    port map (
            in0 => \N__5024\,
            in1 => \N__4455\,
            in2 => \N__4805\,
            in3 => \N__4086\,
            lcout => \sevsegr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_Switch_3_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6556\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \r_SwitchZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7103\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alogicunit.m26_l_fx_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__5357\,
            in1 => \_gnd_net_\,
            in2 => \N__4177\,
            in3 => \_gnd_net_\,
            lcout => \alogicunit.m26_l_fxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sevsegl_RNO_0_1_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__4085\,
            in1 => \N__4789\,
            in2 => \N__4461\,
            in3 => \N__5025\,
            lcout => \sevsegl_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sevsegl_RNO_0_3_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__4790\,
            in1 => \N__5315\,
            in2 => \N__4238\,
            in3 => \N__5130\,
            lcout => \sevsegl_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alogicunit.m26_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__5102\,
            in1 => \N__5018\,
            in2 => \N__5225\,
            in3 => \N__5296\,
            lcout => \alogicunit.result24\,
            ltout => \alogicunit.result24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alogicunit.un1_a_1_cry_3_c_inv_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__4129\,
            in1 => \_gnd_net_\,
            in2 => \N__4137\,
            in3 => \_gnd_net_\,
            lcout => \alogicunit.un1_a_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alogicunit.result_13_iv_5_56_i_o4_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__5209\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5022\,
            lcout => \alogicunit.N_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cu1.track_RNIVBP9_1_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5107\,
            in1 => \N__5301\,
            in2 => \_gnd_net_\,
            in3 => \N__5208\,
            lcout => cu1_track_ns_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cu1.track_RNI9MAL_1_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100111110"
        )
    port map (
            in0 => \N__5207\,
            in1 => \N__5106\,
            in2 => \N__5323\,
            in3 => \N__5020\,
            lcout => \N_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alogicunit.m17_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000001010"
        )
    port map (
            in0 => \N__5021\,
            in1 => \N__5297\,
            in2 => \N__5133\,
            in3 => \N__5210\,
            lcout => \alogicunit.N_41\,
            ltout => \alogicunit.N_41_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alogicunit.result_13_iv_2_182_i_o4_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__5303\,
            in1 => \N__5111\,
            in2 => \N__4494\,
            in3 => \N__5023\,
            lcout => \alogicunit.N_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cu1.track_RNI9MAL_0_1_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010111110"
        )
    port map (
            in0 => \N__5019\,
            in1 => \N__5302\,
            in2 => \N__5132\,
            in3 => \N__5206\,
            lcout => \track_RNI9MAL_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_Count_e_0_2_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__4453\,
            in1 => \N__4321\,
            in2 => \_gnd_net_\,
            in3 => \N__4384\,
            lcout => \r_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7111\,
            ce => \N__4629\,
            sr => \_gnd_net_\
        );

    \Instance2.r_State_RNO_3_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5735\,
            in1 => \N__5504\,
            in2 => \N__5715\,
            in3 => \N__5568\,
            lcout => OPEN,
            ltout => \Instance2.r_Count13_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance2.r_State_RNO_0_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__5543\,
            in1 => \N__6170\,
            in2 => \N__4281\,
            in3 => \N__4635\,
            lcout => \Instance2.r_Count13_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance2.r_Count_RNIIPVO_4_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__5567\,
            in1 => \N__5542\,
            in2 => \N__5505\,
            in3 => \N__5524\,
            lcout => OPEN,
            ltout => \Instance2.un1_r_Count_10lt11_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance2.r_Count_RNINRGT2_12_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100010001"
        )
    port map (
            in0 => \N__5734\,
            in1 => \N__5710\,
            in2 => \N__4278\,
            in3 => \N__4668\,
            lcout => \Instance2.un1_r_Count_10lt17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance2.r_State_RNO_1_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4653\,
            in1 => \N__5759\,
            in2 => \N__4662\,
            in3 => \N__5783\,
            lcout => OPEN,
            ltout => \Instance2.r_Count13_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance2.r_State_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__4871\,
            in1 => \N__4677\,
            in2 => \N__4671\,
            in3 => \N__4916\,
            lcout => \w_Switch_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7099\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance2.r_Count_RNIGGG81_8_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5784\,
            in1 => \N__5479\,
            in2 => \N__5760\,
            in3 => \N__5800\,
            lcout => \Instance2.un1_r_Count_10lto11_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance2.r_State_RNO_5_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__5646\,
            in1 => \N__5525\,
            in2 => \N__5670\,
            in3 => \N__5480\,
            lcout => \Instance2.r_Count13_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance2.r_State_RNO_4_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5801\,
            in1 => \N__5589\,
            in2 => \N__6143\,
            in3 => \N__5603\,
            lcout => \Instance2.r_Count13_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alogicunit.result_13_iv_6_14_i_o4_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__5227\,
            in1 => \N__5145\,
            in2 => \N__5335\,
            in3 => \N__5040\,
            lcout => \alogicunit.N_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance2.r_State_RNO_2_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5692\,
            in2 => \_gnd_net_\,
            in3 => \N__6188\,
            lcout => \Instance2.r_Count13_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance2.r_Count_RNIMF1O1_17_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5641\,
            in1 => \N__6187\,
            in2 => \N__5694\,
            in3 => \N__5665\,
            lcout => \Instance2.un1_r_Count_10lto17_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \click1_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__4760\,
            in1 => \N__4963\,
            in2 => \_gnd_net_\,
            in3 => \N__4625\,
            lcout => \clickZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7104\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alogicunit.result_13_iv_4_98_i_o4_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100100110"
        )
    port map (
            in0 => \N__5226\,
            in1 => \N__5142\,
            in2 => \N__5336\,
            in3 => \N__5037\,
            lcout => \alogicunit.N_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_Switch_2_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4902\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \r_SwitchZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7104\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_Switch_4_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6237\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \r_SwitchZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7104\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance3.r_State_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__6795\,
            in1 => \N__6486\,
            in2 => \N__6537\,
            in3 => \N__6560\,
            lcout => \w_Switch_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7104\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance2.r_State_RNIR73L_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4901\,
            in2 => \_gnd_net_\,
            in3 => \N__4829\,
            lcout => OPEN,
            ltout => \Instance2.click14_sn_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance2.r_State_RNINFUP1_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001101"
        )
    port map (
            in0 => \N__4818\,
            in1 => \N__6236\,
            in2 => \N__4812\,
            in3 => \N__4781\,
            lcout => \Instance2_un1_click13_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alogicunit.result_4_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__4685\,
            in1 => \N__4724\,
            in2 => \_gnd_net_\,
            in3 => \N__4746\,
            lcout => left_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7108\,
            ce => \N__5400\,
            sr => \_gnd_net_\
        );

    \alogicunit.result_6_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__4725\,
            in1 => \N__4686\,
            in2 => \_gnd_net_\,
            in3 => \N__4716\,
            lcout => left_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7108\,
            ce => \N__5400\,
            sr => \_gnd_net_\
        );

    \alogicunit.un1_a_1_cry_1_c_inv_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__6098\,
            in1 => \N__4698\,
            in2 => \_gnd_net_\,
            in3 => \N__5355\,
            lcout => \alogicunit.un1_a_1_cry_1_c_invZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alogicunit.result_13_iv_2_182_i_a2_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110011"
        )
    port map (
            in0 => \N__4990\,
            in1 => \N__5101\,
            in2 => \_gnd_net_\,
            in3 => \N__5201\,
            lcout => \alogicunit.N_102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cu1.track_0_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001100110"
        )
    port map (
            in0 => \N__4955\,
            in1 => \N__5295\,
            in2 => \_gnd_net_\,
            in3 => \N__4991\,
            lcout => current_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cu1.track_1_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__4959\,
            in1 => \N__5320\,
            in2 => \_gnd_net_\,
            in3 => \N__5202\,
            lcout => current_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cu1.track_2_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__5321\,
            in1 => \N__5223\,
            in2 => \N__4964\,
            in3 => \N__5118\,
            lcout => current_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SegInst1.r_HexEncode_i_4_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000010100100"
        )
    port map (
            in0 => \N__6078\,
            in1 => \N__6031\,
            in2 => \N__5989\,
            in3 => \N__5927\,
            lcout => \r_HexEncode_i_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alogicunit.m34_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010111"
        )
    port map (
            in0 => \N__4989\,
            in1 => \N__5319\,
            in2 => \N__5141\,
            in3 => \N__5200\,
            lcout => \alogicunit.N_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \alogicunit.result24_i_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__5100\,
            in1 => \N__4988\,
            in2 => \N__5224\,
            in3 => \N__5294\,
            lcout => \alogicunit.result24_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cu1.track_e_0_3_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5322\,
            in1 => \N__5222\,
            in2 => \_gnd_net_\,
            in3 => \N__5131\,
            lcout => current_state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7115\,
            ce => \N__4965\,
            sr => \_gnd_net_\
        );

    \Instance2.r_State_RNI4PC15_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001111101011"
        )
    port map (
            in0 => \N__4926\,
            in1 => \N__4915\,
            in2 => \N__4878\,
            in3 => \N__4848\,
            lcout => \Instance2.r_Count12_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance4.r_Count_1_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__6455\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5883\,
            lcout => \Instance4.r_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7101\,
            ce => 'H',
            sr => \N__5619\
        );

    \Instance4.r_Count_0_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6454\,
            lcout => \Instance4.r_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7101\,
            ce => 'H',
            sr => \N__5619\
        );

    \Instance4.r_Count_2_cry_1_c_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5882\,
            in2 => \N__6456\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_7_0_\,
            carryout => \Instance4.r_Count_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance4.r_Count_2_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5865\,
            in2 => \_gnd_net_\,
            in3 => \N__5436\,
            lcout => \Instance4.r_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \Instance4.r_Count_2_cry_1\,
            carryout => \Instance4.r_Count_2_cry_2\,
            clk => \N__7095\,
            ce => 'H',
            sr => \N__5620\
        );

    \Instance4.r_Count_3_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5852\,
            in2 => \_gnd_net_\,
            in3 => \N__5433\,
            lcout => \Instance4.r_CountZ0Z_3\,
            ltout => OPEN,
            carryin => \Instance4.r_Count_2_cry_2\,
            carryout => \Instance4.r_Count_2_cry_3\,
            clk => \N__7095\,
            ce => 'H',
            sr => \N__5620\
        );

    \Instance4.r_Count_4_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5838\,
            in2 => \_gnd_net_\,
            in3 => \N__5430\,
            lcout => \Instance4.r_CountZ0Z_4\,
            ltout => OPEN,
            carryin => \Instance4.r_Count_2_cry_3\,
            carryout => \Instance4.r_Count_2_cry_4\,
            clk => \N__7095\,
            ce => 'H',
            sr => \N__5620\
        );

    \Instance4.r_Count_5_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6427\,
            in2 => \_gnd_net_\,
            in3 => \N__5427\,
            lcout => \Instance4.r_CountZ0Z_5\,
            ltout => OPEN,
            carryin => \Instance4.r_Count_2_cry_4\,
            carryout => \Instance4.r_Count_2_cry_5\,
            clk => \N__7095\,
            ce => 'H',
            sr => \N__5620\
        );

    \Instance4.r_Count_6_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6594\,
            in2 => \_gnd_net_\,
            in3 => \N__5424\,
            lcout => \Instance4.r_CountZ0Z_6\,
            ltout => OPEN,
            carryin => \Instance4.r_Count_2_cry_5\,
            carryout => \Instance4.r_Count_2_cry_6\,
            clk => \N__7095\,
            ce => 'H',
            sr => \N__5620\
        );

    \Instance4.r_Count_7_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5819\,
            in2 => \_gnd_net_\,
            in3 => \N__5421\,
            lcout => \Instance4.r_CountZ0Z_7\,
            ltout => OPEN,
            carryin => \Instance4.r_Count_2_cry_6\,
            carryout => \Instance4.r_Count_2_cry_7\,
            clk => \N__7095\,
            ce => 'H',
            sr => \N__5620\
        );

    \Instance4.r_Count_8_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6647\,
            in2 => \_gnd_net_\,
            in3 => \N__5418\,
            lcout => \Instance4.r_CountZ0Z_8\,
            ltout => OPEN,
            carryin => \Instance4.r_Count_2_cry_7\,
            carryout => \Instance4.r_Count_2_cry_8\,
            clk => \N__7095\,
            ce => 'H',
            sr => \N__5620\
        );

    \Instance4.r_Count_9_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6318\,
            in2 => \_gnd_net_\,
            in3 => \N__5463\,
            lcout => \Instance4.r_CountZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_6_8_0_\,
            carryout => \Instance4.r_Count_2_cry_9\,
            clk => \N__7087\,
            ce => 'H',
            sr => \N__5621\
        );

    \Instance4.r_Count_10_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6335\,
            in2 => \_gnd_net_\,
            in3 => \N__5460\,
            lcout => \Instance4.r_CountZ0Z_10\,
            ltout => OPEN,
            carryin => \Instance4.r_Count_2_cry_9\,
            carryout => \Instance4.r_Count_2_cry_10\,
            clk => \N__7087\,
            ce => 'H',
            sr => \N__5621\
        );

    \Instance4.r_Count_11_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6351\,
            in2 => \_gnd_net_\,
            in3 => \N__5457\,
            lcout => \Instance4.r_CountZ0Z_11\,
            ltout => OPEN,
            carryin => \Instance4.r_Count_2_cry_10\,
            carryout => \Instance4.r_Count_2_cry_11\,
            clk => \N__7087\,
            ce => 'H',
            sr => \N__5621\
        );

    \Instance4.r_Count_12_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6282\,
            in2 => \_gnd_net_\,
            in3 => \N__5454\,
            lcout => \Instance4.r_CountZ0Z_12\,
            ltout => OPEN,
            carryin => \Instance4.r_Count_2_cry_11\,
            carryout => \Instance4.r_Count_2_cry_12\,
            clk => \N__7087\,
            ce => 'H',
            sr => \N__5621\
        );

    \Instance4.r_Count_13_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6300\,
            in2 => \_gnd_net_\,
            in3 => \N__5451\,
            lcout => \Instance4.r_CountZ0Z_13\,
            ltout => OPEN,
            carryin => \Instance4.r_Count_2_cry_12\,
            carryout => \Instance4.r_Count_2_cry_13\,
            clk => \N__7087\,
            ce => 'H',
            sr => \N__5621\
        );

    \Instance4.r_Count_14_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6389\,
            in2 => \_gnd_net_\,
            in3 => \N__5448\,
            lcout => \Instance4.r_CountZ0Z_14\,
            ltout => OPEN,
            carryin => \Instance4.r_Count_2_cry_13\,
            carryout => \Instance4.r_Count_2_cry_14\,
            clk => \N__7087\,
            ce => 'H',
            sr => \N__5621\
        );

    \Instance4.r_Count_15_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6630\,
            in2 => \_gnd_net_\,
            in3 => \N__5445\,
            lcout => \Instance4.r_CountZ0Z_15\,
            ltout => OPEN,
            carryin => \Instance4.r_Count_2_cry_14\,
            carryout => \Instance4.r_Count_2_cry_15\,
            clk => \N__7087\,
            ce => 'H',
            sr => \N__5621\
        );

    \Instance4.r_Count_16_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6611\,
            in2 => \_gnd_net_\,
            in3 => \N__5442\,
            lcout => \Instance4.r_CountZ0Z_16\,
            ltout => OPEN,
            carryin => \Instance4.r_Count_2_cry_15\,
            carryout => \Instance4.r_Count_2_cry_16\,
            clk => \N__7087\,
            ce => 'H',
            sr => \N__5621\
        );

    \Instance4.r_Count_17_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6372\,
            in2 => \_gnd_net_\,
            in3 => \N__5439\,
            lcout => \Instance4.r_CountZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7096\,
            ce => 'H',
            sr => \N__5622\
        );

    \Instance2.r_Count_2_cry_1_c_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6144\,
            in2 => \N__6171\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_10_0_\,
            carryout => \Instance2.r_Count_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance2.r_Count_2_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5604\,
            in2 => \_gnd_net_\,
            in3 => \N__5592\,
            lcout => \Instance2.r_Count_0_2\,
            ltout => OPEN,
            carryin => \Instance2.r_Count_2_cry_1\,
            carryout => \Instance2.r_Count_2_cry_2\,
            clk => \N__7100\,
            ce => 'H',
            sr => \N__6120\
        );

    \Instance2.r_Count_3_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5582\,
            in2 => \_gnd_net_\,
            in3 => \N__5571\,
            lcout => \Instance2.r_Count_0_3\,
            ltout => OPEN,
            carryin => \Instance2.r_Count_2_cry_2\,
            carryout => \Instance2.r_Count_2_cry_3\,
            clk => \N__7100\,
            ce => 'H',
            sr => \N__6120\
        );

    \Instance2.r_Count_4_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5566\,
            in2 => \_gnd_net_\,
            in3 => \N__5547\,
            lcout => \Instance2.r_CountZ0Z_4\,
            ltout => OPEN,
            carryin => \Instance2.r_Count_2_cry_3\,
            carryout => \Instance2.r_Count_2_cry_4\,
            clk => \N__7100\,
            ce => 'H',
            sr => \N__6120\
        );

    \Instance2.r_Count_5_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5544\,
            in2 => \_gnd_net_\,
            in3 => \N__5529\,
            lcout => \Instance2.r_CountZ0Z_5\,
            ltout => OPEN,
            carryin => \Instance2.r_Count_2_cry_4\,
            carryout => \Instance2.r_Count_2_cry_5\,
            clk => \N__7100\,
            ce => 'H',
            sr => \N__6120\
        );

    \Instance2.r_Count_6_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5526\,
            in2 => \_gnd_net_\,
            in3 => \N__5508\,
            lcout => \Instance2.r_CountZ0Z_6\,
            ltout => OPEN,
            carryin => \Instance2.r_Count_2_cry_5\,
            carryout => \Instance2.r_Count_2_cry_6\,
            clk => \N__7100\,
            ce => 'H',
            sr => \N__6120\
        );

    \Instance2.r_Count_7_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5503\,
            in2 => \_gnd_net_\,
            in3 => \N__5484\,
            lcout => \Instance2.r_CountZ0Z_7\,
            ltout => OPEN,
            carryin => \Instance2.r_Count_2_cry_6\,
            carryout => \Instance2.r_Count_2_cry_7\,
            clk => \N__7100\,
            ce => 'H',
            sr => \N__6120\
        );

    \Instance2.r_Count_8_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5481\,
            in2 => \_gnd_net_\,
            in3 => \N__5466\,
            lcout => \Instance2.r_CountZ0Z_8\,
            ltout => OPEN,
            carryin => \Instance2.r_Count_2_cry_7\,
            carryout => \Instance2.r_Count_2_cry_8\,
            clk => \N__7100\,
            ce => 'H',
            sr => \N__6120\
        );

    \Instance2.r_Count_9_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5802\,
            in2 => \_gnd_net_\,
            in3 => \N__5787\,
            lcout => \Instance2.r_CountZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_6_11_0_\,
            carryout => \Instance2.r_Count_2_cry_9\,
            clk => \N__7105\,
            ce => 'H',
            sr => \N__6119\
        );

    \Instance2.r_Count_10_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5782\,
            in2 => \_gnd_net_\,
            in3 => \N__5763\,
            lcout => \Instance2.r_CountZ0Z_10\,
            ltout => OPEN,
            carryin => \Instance2.r_Count_2_cry_9\,
            carryout => \Instance2.r_Count_2_cry_10\,
            clk => \N__7105\,
            ce => 'H',
            sr => \N__6119\
        );

    \Instance2.r_Count_11_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5758\,
            in2 => \_gnd_net_\,
            in3 => \N__5739\,
            lcout => \Instance2.r_CountZ0Z_11\,
            ltout => OPEN,
            carryin => \Instance2.r_Count_2_cry_10\,
            carryout => \Instance2.r_Count_2_cry_11\,
            clk => \N__7105\,
            ce => 'H',
            sr => \N__6119\
        );

    \Instance2.r_Count_12_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5736\,
            in2 => \_gnd_net_\,
            in3 => \N__5718\,
            lcout => \Instance2.r_CountZ0Z_12\,
            ltout => OPEN,
            carryin => \Instance2.r_Count_2_cry_11\,
            carryout => \Instance2.r_Count_2_cry_12\,
            clk => \N__7105\,
            ce => 'H',
            sr => \N__6119\
        );

    \Instance2.r_Count_13_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5714\,
            in2 => \_gnd_net_\,
            in3 => \N__5697\,
            lcout => \Instance2.r_CountZ0Z_13\,
            ltout => OPEN,
            carryin => \Instance2.r_Count_2_cry_12\,
            carryout => \Instance2.r_Count_2_cry_13\,
            clk => \N__7105\,
            ce => 'H',
            sr => \N__6119\
        );

    \Instance2.r_Count_14_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5693\,
            in2 => \_gnd_net_\,
            in3 => \N__5673\,
            lcout => \Instance2.r_CountZ0Z_14\,
            ltout => OPEN,
            carryin => \Instance2.r_Count_2_cry_13\,
            carryout => \Instance2.r_Count_2_cry_14\,
            clk => \N__7105\,
            ce => 'H',
            sr => \N__6119\
        );

    \Instance2.r_Count_15_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5669\,
            in2 => \_gnd_net_\,
            in3 => \N__5649\,
            lcout => \Instance2.r_CountZ0Z_15\,
            ltout => OPEN,
            carryin => \Instance2.r_Count_2_cry_14\,
            carryout => \Instance2.r_Count_2_cry_15\,
            clk => \N__7105\,
            ce => 'H',
            sr => \N__6119\
        );

    \Instance2.r_Count_16_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5645\,
            in2 => \_gnd_net_\,
            in3 => \N__5625\,
            lcout => \Instance2.r_CountZ0Z_16\,
            ltout => OPEN,
            carryin => \Instance2.r_Count_2_cry_15\,
            carryout => \Instance2.r_Count_2_cry_16\,
            clk => \N__7105\,
            ce => 'H',
            sr => \N__6119\
        );

    \Instance2.r_Count_17_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6189\,
            in2 => \_gnd_net_\,
            in3 => \N__6192\,
            lcout => \Instance2.r_CountZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7109\,
            ce => 'H',
            sr => \N__6118\
        );

    \Instance2.r_Count_0_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6165\,
            lcout => \Instance2.r_Count_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7109\,
            ce => 'H',
            sr => \N__6118\
        );

    \Instance2.r_Count_1_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__6166\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6142\,
            lcout => \Instance2.r_Count_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7109\,
            ce => 'H',
            sr => \N__6118\
        );

    \CONSTANT_ONE_LUT4_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SegInst1.r_HexEncode_i_3_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100101000010"
        )
    port map (
            in0 => \N__6077\,
            in1 => \N__6033\,
            in2 => \N__5991\,
            in3 => \N__5934\,
            lcout => \r_HexEncode_i_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7116\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SegInst1.r_HexEncode_i_2_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001111100000010"
        )
    port map (
            in0 => \N__6076\,
            in1 => \N__6032\,
            in2 => \N__5990\,
            in3 => \N__5933\,
            lcout => \r_HexEncode_i_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7116\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance4.r_State_RNO_4_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5881\,
            in1 => \N__5864\,
            in2 => \N__5853\,
            in3 => \N__6317\,
            lcout => \Instance4.r_Count13_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance4.r_Count_RNIQHQE_4_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__5818\,
            in1 => \N__5836\,
            in2 => \N__6429\,
            in3 => \N__6592\,
            lcout => \Instance4.un1_r_Count_10lt11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance4.r_State_RNO_3_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5837\,
            in1 => \N__6299\,
            in2 => \N__5823\,
            in3 => \N__6281\,
            lcout => OPEN,
            ltout => \Instance4.r_Count13_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance4.r_State_RNO_0_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__6357\,
            in1 => \N__6453\,
            in2 => \N__6432\,
            in3 => \N__6428\,
            lcout => \Instance4.r_Count13_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance4.r_State_RNO_1_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6334\,
            in1 => \N__6408\,
            in2 => \N__6576\,
            in3 => \N__6350\,
            lcout => OPEN,
            ltout => \Instance4.r_Count13_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance4.r_State_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__6227\,
            in1 => \N__6254\,
            in2 => \N__6402\,
            in3 => \N__6399\,
            lcout => \w_Switch_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7091\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance4.r_Count_RNIUFK81_17_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6370\,
            in1 => \N__6628\,
            in2 => \N__6390\,
            in3 => \N__6607\,
            lcout => \Instance4.un1_r_Count_10lto17_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance4.r_State_RNO_2_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6388\,
            in2 => \_gnd_net_\,
            in3 => \N__6371\,
            lcout => \Instance4.r_Count13_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance4.r_Count_RNIOCNR_8_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6646\,
            in1 => \N__6349\,
            in2 => \N__6336\,
            in3 => \N__6316\,
            lcout => OPEN,
            ltout => \Instance4.un1_r_Count_10lto11_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance4.r_Count_RNIB0SU1_12_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010001"
        )
    port map (
            in0 => \N__6298\,
            in1 => \N__6280\,
            in2 => \N__6264\,
            in3 => \N__6261\,
            lcout => OPEN,
            ltout => \Instance4.un1_r_Count_10lt17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance4.r_State_RNI4ONP3_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111110011001"
        )
    port map (
            in0 => \N__6255\,
            in1 => \N__6226\,
            in2 => \N__6213\,
            in3 => \N__6210\,
            lcout => \Instance4.r_Count12_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance4.r_State_RNO_5_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6648\,
            in1 => \N__6629\,
            in2 => \N__6612\,
            in3 => \N__6593\,
            lcout => \Instance4.r_Count13_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance3.r_Count_RNI1E6U3_12_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100000011"
        )
    port map (
            in0 => \N__6474\,
            in1 => \N__6814\,
            in2 => \N__6846\,
            in3 => \N__6468\,
            lcout => OPEN,
            ltout => \Instance3.un1_r_Count_10lt17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance3.r_State_RNIK8IT5_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111110011001"
        )
    port map (
            in0 => \N__6567\,
            in1 => \N__6530\,
            in2 => \N__6501\,
            in3 => \N__6777\,
            lcout => \Instance3.r_Count12_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance3.r_State_RNO_3_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6841\,
            in1 => \N__6956\,
            in2 => \N__6819\,
            in3 => \N__6686\,
            lcout => OPEN,
            ltout => \Instance3.r_Count13_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance3.r_State_RNO_0_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__6668\,
            in1 => \N__7167\,
            in2 => \N__6489\,
            in3 => \N__6462\,
            lcout => \Instance3.r_Count13_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance3.r_Count_RNIM5TJ1_4_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__6669\,
            in1 => \N__6685\,
            in2 => \N__6981\,
            in3 => \N__6955\,
            lcout => \Instance3.un1_r_Count_10lt11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance3.r_Count_RNIKU3I1_10_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6870\,
            in1 => \N__6937\,
            in2 => \N__6897\,
            in3 => \N__6916\,
            lcout => \Instance3.un1_r_Count_10lto11_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance3.r_State_RNO_2_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7249\,
            in2 => \_gnd_net_\,
            in3 => \N__7181\,
            lcout => \Instance3.r_Count13_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance3.r_State_RNO_4_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6719\,
            in1 => \N__7137\,
            in2 => \N__6705\,
            in3 => \N__6917\,
            lcout => OPEN,
            ltout => \Instance3.r_Count13_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance3.r_State_RNO_1_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__6783\,
            in1 => \N__6868\,
            in2 => \N__6798\,
            in3 => \N__6892\,
            lcout => \Instance3.r_Count13_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance3.r_State_RNO_5_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__7205\,
            in1 => \N__6979\,
            in2 => \N__7230\,
            in3 => \N__6938\,
            lcout => \Instance3.r_Count13_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance3.r_Count_RNIQVAG1_17_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7180\,
            in1 => \N__7225\,
            in2 => \N__7251\,
            in3 => \N__7204\,
            lcout => \Instance3.un1_r_Count_10lto17_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_1_1_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6771\,
            lcout => \o_LED_1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance3.r_Count_2_cry_1_c_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7135\,
            in2 => \N__7163\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => \Instance3.r_Count_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Instance3.r_Count_2_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6720\,
            in2 => \_gnd_net_\,
            in3 => \N__6708\,
            lcout => \Instance3.r_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \Instance3.r_Count_2_cry_1\,
            carryout => \Instance3.r_Count_2_cry_2\,
            clk => \N__7106\,
            ce => 'H',
            sr => \N__6999\
        );

    \Instance3.r_Count_3_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6704\,
            in2 => \_gnd_net_\,
            in3 => \N__6690\,
            lcout => \Instance3.r_CountZ0Z_3\,
            ltout => OPEN,
            carryin => \Instance3.r_Count_2_cry_2\,
            carryout => \Instance3.r_Count_2_cry_3\,
            clk => \N__7106\,
            ce => 'H',
            sr => \N__6999\
        );

    \Instance3.r_Count_4_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6687\,
            in2 => \_gnd_net_\,
            in3 => \N__6672\,
            lcout => \Instance3.r_CountZ0Z_4\,
            ltout => OPEN,
            carryin => \Instance3.r_Count_2_cry_3\,
            carryout => \Instance3.r_Count_2_cry_4\,
            clk => \N__7106\,
            ce => 'H',
            sr => \N__6999\
        );

    \Instance3.r_Count_5_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6667\,
            in2 => \_gnd_net_\,
            in3 => \N__6984\,
            lcout => \Instance3.r_CountZ0Z_5\,
            ltout => OPEN,
            carryin => \Instance3.r_Count_2_cry_4\,
            carryout => \Instance3.r_Count_2_cry_5\,
            clk => \N__7106\,
            ce => 'H',
            sr => \N__6999\
        );

    \Instance3.r_Count_6_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6980\,
            in2 => \_gnd_net_\,
            in3 => \N__6960\,
            lcout => \Instance3.r_CountZ0Z_6\,
            ltout => OPEN,
            carryin => \Instance3.r_Count_2_cry_5\,
            carryout => \Instance3.r_Count_2_cry_6\,
            clk => \N__7106\,
            ce => 'H',
            sr => \N__6999\
        );

    \Instance3.r_Count_7_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6957\,
            in2 => \_gnd_net_\,
            in3 => \N__6942\,
            lcout => \Instance3.r_CountZ0Z_7\,
            ltout => OPEN,
            carryin => \Instance3.r_Count_2_cry_6\,
            carryout => \Instance3.r_Count_2_cry_7\,
            clk => \N__7106\,
            ce => 'H',
            sr => \N__6999\
        );

    \Instance3.r_Count_8_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6939\,
            in2 => \_gnd_net_\,
            in3 => \N__6921\,
            lcout => \Instance3.r_CountZ0Z_8\,
            ltout => OPEN,
            carryin => \Instance3.r_Count_2_cry_7\,
            carryout => \Instance3.r_Count_2_cry_8\,
            clk => \N__7106\,
            ce => 'H',
            sr => \N__6999\
        );

    \Instance3.r_Count_9_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6918\,
            in2 => \_gnd_net_\,
            in3 => \N__6900\,
            lcout => \Instance3.r_CountZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => \Instance3.r_Count_2_cry_9\,
            clk => \N__7110\,
            ce => 'H',
            sr => \N__7001\
        );

    \Instance3.r_Count_10_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6893\,
            in2 => \_gnd_net_\,
            in3 => \N__6873\,
            lcout => \Instance3.r_CountZ0Z_10\,
            ltout => OPEN,
            carryin => \Instance3.r_Count_2_cry_9\,
            carryout => \Instance3.r_Count_2_cry_10\,
            clk => \N__7110\,
            ce => 'H',
            sr => \N__7001\
        );

    \Instance3.r_Count_11_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6869\,
            in2 => \_gnd_net_\,
            in3 => \N__6849\,
            lcout => \Instance3.r_CountZ0Z_11\,
            ltout => OPEN,
            carryin => \Instance3.r_Count_2_cry_10\,
            carryout => \Instance3.r_Count_2_cry_11\,
            clk => \N__7110\,
            ce => 'H',
            sr => \N__7001\
        );

    \Instance3.r_Count_12_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6842\,
            in2 => \_gnd_net_\,
            in3 => \N__6822\,
            lcout => \Instance3.r_CountZ0Z_12\,
            ltout => OPEN,
            carryin => \Instance3.r_Count_2_cry_11\,
            carryout => \Instance3.r_Count_2_cry_12\,
            clk => \N__7110\,
            ce => 'H',
            sr => \N__7001\
        );

    \Instance3.r_Count_13_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6818\,
            in2 => \_gnd_net_\,
            in3 => \N__6801\,
            lcout => \Instance3.r_CountZ0Z_13\,
            ltout => OPEN,
            carryin => \Instance3.r_Count_2_cry_12\,
            carryout => \Instance3.r_Count_2_cry_13\,
            clk => \N__7110\,
            ce => 'H',
            sr => \N__7001\
        );

    \Instance3.r_Count_14_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7250\,
            in2 => \_gnd_net_\,
            in3 => \N__7233\,
            lcout => \Instance3.r_CountZ0Z_14\,
            ltout => OPEN,
            carryin => \Instance3.r_Count_2_cry_13\,
            carryout => \Instance3.r_Count_2_cry_14\,
            clk => \N__7110\,
            ce => 'H',
            sr => \N__7001\
        );

    \Instance3.r_Count_15_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7229\,
            in2 => \_gnd_net_\,
            in3 => \N__7209\,
            lcout => \Instance3.r_CountZ0Z_15\,
            ltout => OPEN,
            carryin => \Instance3.r_Count_2_cry_14\,
            carryout => \Instance3.r_Count_2_cry_15\,
            clk => \N__7110\,
            ce => 'H',
            sr => \N__7001\
        );

    \Instance3.r_Count_16_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7206\,
            in2 => \_gnd_net_\,
            in3 => \N__7188\,
            lcout => \Instance3.r_CountZ0Z_16\,
            ltout => OPEN,
            carryin => \Instance3.r_Count_2_cry_15\,
            carryout => \Instance3.r_Count_2_cry_16\,
            clk => \N__7110\,
            ce => 'H',
            sr => \N__7001\
        );

    \Instance3.r_Count_17_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7182\,
            in2 => \_gnd_net_\,
            in3 => \N__7185\,
            lcout => \Instance3.r_CountZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7113\,
            ce => 'H',
            sr => \N__7002\
        );

    \Instance3.r_Count_0_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7161\,
            lcout => \Instance3.r_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7114\,
            ce => 'H',
            sr => \N__7000\
        );

    \Instance3.r_Count_1_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__7162\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7136\,
            lcout => \Instance3.r_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7114\,
            ce => 'H',
            sr => \N__7000\
        );
end \INTERFACE\;
