// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Aug 6 2023 18:36:21

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "simpleprocessor_top" view "INTERFACE"

module simpleprocessor_top (
    o_Segment2_F,
    o_Segment1_D,
    o_LED_1,
    o_Segment2_A,
    o_Segment1_E,
    o_Segment2_D,
    o_Segment1_F,
    o_Segment1_B,
    o_LED_3,
    i_Switch_4,
    i_Clk,
    o_Segment2_G,
    o_Segment2_C,
    o_Segment1_G,
    o_Segment1_C,
    o_LED_2,
    i_Switch_1,
    o_Segment2_B,
    i_Switch_2,
    o_Segment2_E,
    o_Segment1_A,
    o_LED_4,
    i_Switch_3);

    output o_Segment2_F;
    output o_Segment1_D;
    output o_LED_1;
    output o_Segment2_A;
    output o_Segment1_E;
    output o_Segment2_D;
    output o_Segment1_F;
    output o_Segment1_B;
    output o_LED_3;
    input i_Switch_4;
    input i_Clk;
    output o_Segment2_G;
    output o_Segment2_C;
    output o_Segment1_G;
    output o_Segment1_C;
    output o_LED_2;
    input i_Switch_1;
    output o_Segment2_B;
    input i_Switch_2;
    output o_Segment2_E;
    output o_Segment1_A;
    output o_LED_4;
    input i_Switch_3;

    wire N__7470;
    wire N__7469;
    wire N__7468;
    wire N__7459;
    wire N__7458;
    wire N__7457;
    wire N__7450;
    wire N__7449;
    wire N__7448;
    wire N__7441;
    wire N__7440;
    wire N__7439;
    wire N__7432;
    wire N__7431;
    wire N__7430;
    wire N__7423;
    wire N__7422;
    wire N__7421;
    wire N__7414;
    wire N__7413;
    wire N__7412;
    wire N__7405;
    wire N__7404;
    wire N__7403;
    wire N__7396;
    wire N__7395;
    wire N__7394;
    wire N__7387;
    wire N__7386;
    wire N__7385;
    wire N__7378;
    wire N__7377;
    wire N__7376;
    wire N__7369;
    wire N__7368;
    wire N__7367;
    wire N__7360;
    wire N__7359;
    wire N__7358;
    wire N__7351;
    wire N__7350;
    wire N__7349;
    wire N__7342;
    wire N__7341;
    wire N__7340;
    wire N__7333;
    wire N__7332;
    wire N__7331;
    wire N__7324;
    wire N__7323;
    wire N__7322;
    wire N__7315;
    wire N__7314;
    wire N__7313;
    wire N__7306;
    wire N__7305;
    wire N__7304;
    wire N__7297;
    wire N__7296;
    wire N__7295;
    wire N__7288;
    wire N__7287;
    wire N__7286;
    wire N__7279;
    wire N__7278;
    wire N__7277;
    wire N__7270;
    wire N__7269;
    wire N__7268;
    wire N__7251;
    wire N__7250;
    wire N__7249;
    wire N__7246;
    wire N__7243;
    wire N__7238;
    wire N__7233;
    wire N__7230;
    wire N__7229;
    wire N__7226;
    wire N__7225;
    wire N__7222;
    wire N__7219;
    wire N__7216;
    wire N__7209;
    wire N__7206;
    wire N__7205;
    wire N__7204;
    wire N__7201;
    wire N__7198;
    wire N__7195;
    wire N__7188;
    wire N__7185;
    wire N__7182;
    wire N__7181;
    wire N__7180;
    wire N__7177;
    wire N__7172;
    wire N__7167;
    wire N__7164;
    wire N__7163;
    wire N__7162;
    wire N__7161;
    wire N__7158;
    wire N__7155;
    wire N__7150;
    wire N__7147;
    wire N__7144;
    wire N__7137;
    wire N__7136;
    wire N__7135;
    wire N__7132;
    wire N__7129;
    wire N__7126;
    wire N__7123;
    wire N__7116;
    wire N__7115;
    wire N__7114;
    wire N__7113;
    wire N__7112;
    wire N__7111;
    wire N__7110;
    wire N__7109;
    wire N__7108;
    wire N__7107;
    wire N__7106;
    wire N__7105;
    wire N__7104;
    wire N__7103;
    wire N__7102;
    wire N__7101;
    wire N__7100;
    wire N__7099;
    wire N__7098;
    wire N__7097;
    wire N__7096;
    wire N__7095;
    wire N__7094;
    wire N__7093;
    wire N__7092;
    wire N__7091;
    wire N__7090;
    wire N__7089;
    wire N__7088;
    wire N__7087;
    wire N__7086;
    wire N__7085;
    wire N__7084;
    wire N__7083;
    wire N__7082;
    wire N__7081;
    wire N__7008;
    wire N__7005;
    wire N__7002;
    wire N__7001;
    wire N__7000;
    wire N__6999;
    wire N__6990;
    wire N__6987;
    wire N__6984;
    wire N__6981;
    wire N__6980;
    wire N__6979;
    wire N__6976;
    wire N__6973;
    wire N__6970;
    wire N__6967;
    wire N__6960;
    wire N__6957;
    wire N__6956;
    wire N__6955;
    wire N__6952;
    wire N__6947;
    wire N__6942;
    wire N__6939;
    wire N__6938;
    wire N__6937;
    wire N__6934;
    wire N__6931;
    wire N__6928;
    wire N__6921;
    wire N__6918;
    wire N__6917;
    wire N__6916;
    wire N__6913;
    wire N__6910;
    wire N__6907;
    wire N__6900;
    wire N__6897;
    wire N__6894;
    wire N__6893;
    wire N__6892;
    wire N__6889;
    wire N__6886;
    wire N__6883;
    wire N__6880;
    wire N__6873;
    wire N__6870;
    wire N__6869;
    wire N__6868;
    wire N__6865;
    wire N__6862;
    wire N__6859;
    wire N__6856;
    wire N__6849;
    wire N__6846;
    wire N__6843;
    wire N__6842;
    wire N__6841;
    wire N__6838;
    wire N__6835;
    wire N__6832;
    wire N__6829;
    wire N__6822;
    wire N__6819;
    wire N__6818;
    wire N__6815;
    wire N__6814;
    wire N__6811;
    wire N__6806;
    wire N__6801;
    wire N__6798;
    wire N__6795;
    wire N__6792;
    wire N__6789;
    wire N__6786;
    wire N__6783;
    wire N__6780;
    wire N__6777;
    wire N__6774;
    wire N__6771;
    wire N__6768;
    wire N__6765;
    wire N__6762;
    wire N__6759;
    wire N__6758;
    wire N__6757;
    wire N__6754;
    wire N__6751;
    wire N__6748;
    wire N__6747;
    wire N__6744;
    wire N__6739;
    wire N__6736;
    wire N__6733;
    wire N__6730;
    wire N__6727;
    wire N__6720;
    wire N__6719;
    wire N__6716;
    wire N__6713;
    wire N__6708;
    wire N__6705;
    wire N__6704;
    wire N__6701;
    wire N__6698;
    wire N__6695;
    wire N__6690;
    wire N__6687;
    wire N__6686;
    wire N__6685;
    wire N__6682;
    wire N__6677;
    wire N__6672;
    wire N__6669;
    wire N__6668;
    wire N__6667;
    wire N__6664;
    wire N__6661;
    wire N__6658;
    wire N__6655;
    wire N__6648;
    wire N__6647;
    wire N__6646;
    wire N__6643;
    wire N__6640;
    wire N__6637;
    wire N__6630;
    wire N__6629;
    wire N__6628;
    wire N__6625;
    wire N__6622;
    wire N__6619;
    wire N__6612;
    wire N__6611;
    wire N__6608;
    wire N__6607;
    wire N__6604;
    wire N__6599;
    wire N__6594;
    wire N__6593;
    wire N__6592;
    wire N__6589;
    wire N__6586;
    wire N__6583;
    wire N__6576;
    wire N__6573;
    wire N__6570;
    wire N__6567;
    wire N__6564;
    wire N__6561;
    wire N__6560;
    wire N__6557;
    wire N__6556;
    wire N__6555;
    wire N__6552;
    wire N__6549;
    wire N__6544;
    wire N__6537;
    wire N__6534;
    wire N__6531;
    wire N__6530;
    wire N__6527;
    wire N__6524;
    wire N__6521;
    wire N__6518;
    wire N__6515;
    wire N__6512;
    wire N__6509;
    wire N__6506;
    wire N__6501;
    wire N__6498;
    wire N__6495;
    wire N__6492;
    wire N__6489;
    wire N__6486;
    wire N__6483;
    wire N__6480;
    wire N__6477;
    wire N__6474;
    wire N__6471;
    wire N__6468;
    wire N__6465;
    wire N__6462;
    wire N__6459;
    wire N__6456;
    wire N__6455;
    wire N__6454;
    wire N__6453;
    wire N__6450;
    wire N__6445;
    wire N__6442;
    wire N__6439;
    wire N__6432;
    wire N__6429;
    wire N__6428;
    wire N__6427;
    wire N__6424;
    wire N__6421;
    wire N__6418;
    wire N__6415;
    wire N__6408;
    wire N__6405;
    wire N__6402;
    wire N__6399;
    wire N__6396;
    wire N__6393;
    wire N__6390;
    wire N__6389;
    wire N__6388;
    wire N__6385;
    wire N__6382;
    wire N__6377;
    wire N__6372;
    wire N__6371;
    wire N__6370;
    wire N__6367;
    wire N__6362;
    wire N__6357;
    wire N__6354;
    wire N__6351;
    wire N__6350;
    wire N__6349;
    wire N__6346;
    wire N__6341;
    wire N__6336;
    wire N__6335;
    wire N__6334;
    wire N__6331;
    wire N__6328;
    wire N__6323;
    wire N__6318;
    wire N__6317;
    wire N__6316;
    wire N__6313;
    wire N__6310;
    wire N__6307;
    wire N__6300;
    wire N__6299;
    wire N__6298;
    wire N__6295;
    wire N__6292;
    wire N__6289;
    wire N__6282;
    wire N__6281;
    wire N__6280;
    wire N__6277;
    wire N__6274;
    wire N__6271;
    wire N__6264;
    wire N__6261;
    wire N__6258;
    wire N__6255;
    wire N__6254;
    wire N__6249;
    wire N__6246;
    wire N__6243;
    wire N__6240;
    wire N__6237;
    wire N__6236;
    wire N__6231;
    wire N__6228;
    wire N__6227;
    wire N__6226;
    wire N__6223;
    wire N__6218;
    wire N__6213;
    wire N__6210;
    wire N__6207;
    wire N__6204;
    wire N__6201;
    wire N__6198;
    wire N__6195;
    wire N__6192;
    wire N__6189;
    wire N__6188;
    wire N__6187;
    wire N__6184;
    wire N__6181;
    wire N__6178;
    wire N__6171;
    wire N__6170;
    wire N__6167;
    wire N__6166;
    wire N__6165;
    wire N__6162;
    wire N__6159;
    wire N__6154;
    wire N__6149;
    wire N__6144;
    wire N__6143;
    wire N__6142;
    wire N__6139;
    wire N__6136;
    wire N__6133;
    wire N__6130;
    wire N__6127;
    wire N__6120;
    wire N__6119;
    wire N__6118;
    wire N__6111;
    wire N__6108;
    wire N__6105;
    wire N__6102;
    wire N__6099;
    wire N__6098;
    wire N__6095;
    wire N__6092;
    wire N__6087;
    wire N__6084;
    wire N__6081;
    wire N__6078;
    wire N__6077;
    wire N__6076;
    wire N__6073;
    wire N__6068;
    wire N__6067;
    wire N__6066;
    wire N__6061;
    wire N__6060;
    wire N__6059;
    wire N__6054;
    wire N__6051;
    wire N__6046;
    wire N__6043;
    wire N__6040;
    wire N__6033;
    wire N__6032;
    wire N__6031;
    wire N__6030;
    wire N__6025;
    wire N__6022;
    wire N__6019;
    wire N__6018;
    wire N__6017;
    wire N__6016;
    wire N__6011;
    wire N__6006;
    wire N__6001;
    wire N__5998;
    wire N__5991;
    wire N__5990;
    wire N__5989;
    wire N__5986;
    wire N__5983;
    wire N__5980;
    wire N__5975;
    wire N__5972;
    wire N__5971;
    wire N__5970;
    wire N__5969;
    wire N__5964;
    wire N__5963;
    wire N__5960;
    wire N__5957;
    wire N__5954;
    wire N__5951;
    wire N__5946;
    wire N__5941;
    wire N__5934;
    wire N__5933;
    wire N__5928;
    wire N__5927;
    wire N__5924;
    wire N__5921;
    wire N__5916;
    wire N__5915;
    wire N__5914;
    wire N__5913;
    wire N__5912;
    wire N__5909;
    wire N__5904;
    wire N__5899;
    wire N__5892;
    wire N__5889;
    wire N__5886;
    wire N__5883;
    wire N__5882;
    wire N__5881;
    wire N__5878;
    wire N__5875;
    wire N__5872;
    wire N__5865;
    wire N__5864;
    wire N__5861;
    wire N__5858;
    wire N__5853;
    wire N__5852;
    wire N__5849;
    wire N__5846;
    wire N__5843;
    wire N__5838;
    wire N__5837;
    wire N__5836;
    wire N__5833;
    wire N__5828;
    wire N__5823;
    wire N__5820;
    wire N__5819;
    wire N__5818;
    wire N__5815;
    wire N__5812;
    wire N__5809;
    wire N__5802;
    wire N__5801;
    wire N__5800;
    wire N__5797;
    wire N__5792;
    wire N__5787;
    wire N__5784;
    wire N__5783;
    wire N__5782;
    wire N__5779;
    wire N__5776;
    wire N__5773;
    wire N__5770;
    wire N__5763;
    wire N__5760;
    wire N__5759;
    wire N__5758;
    wire N__5755;
    wire N__5752;
    wire N__5749;
    wire N__5746;
    wire N__5739;
    wire N__5736;
    wire N__5735;
    wire N__5734;
    wire N__5731;
    wire N__5728;
    wire N__5725;
    wire N__5718;
    wire N__5715;
    wire N__5714;
    wire N__5711;
    wire N__5710;
    wire N__5707;
    wire N__5702;
    wire N__5697;
    wire N__5694;
    wire N__5693;
    wire N__5692;
    wire N__5689;
    wire N__5686;
    wire N__5683;
    wire N__5680;
    wire N__5673;
    wire N__5670;
    wire N__5669;
    wire N__5666;
    wire N__5665;
    wire N__5662;
    wire N__5659;
    wire N__5656;
    wire N__5649;
    wire N__5646;
    wire N__5645;
    wire N__5642;
    wire N__5641;
    wire N__5638;
    wire N__5635;
    wire N__5632;
    wire N__5625;
    wire N__5622;
    wire N__5621;
    wire N__5620;
    wire N__5619;
    wire N__5610;
    wire N__5607;
    wire N__5604;
    wire N__5603;
    wire N__5600;
    wire N__5597;
    wire N__5592;
    wire N__5589;
    wire N__5586;
    wire N__5583;
    wire N__5582;
    wire N__5579;
    wire N__5576;
    wire N__5571;
    wire N__5568;
    wire N__5567;
    wire N__5566;
    wire N__5563;
    wire N__5560;
    wire N__5557;
    wire N__5552;
    wire N__5547;
    wire N__5544;
    wire N__5543;
    wire N__5542;
    wire N__5539;
    wire N__5534;
    wire N__5529;
    wire N__5526;
    wire N__5525;
    wire N__5524;
    wire N__5521;
    wire N__5518;
    wire N__5515;
    wire N__5508;
    wire N__5505;
    wire N__5504;
    wire N__5503;
    wire N__5500;
    wire N__5497;
    wire N__5494;
    wire N__5491;
    wire N__5484;
    wire N__5481;
    wire N__5480;
    wire N__5479;
    wire N__5476;
    wire N__5471;
    wire N__5466;
    wire N__5463;
    wire N__5460;
    wire N__5457;
    wire N__5454;
    wire N__5451;
    wire N__5448;
    wire N__5445;
    wire N__5442;
    wire N__5439;
    wire N__5436;
    wire N__5433;
    wire N__5430;
    wire N__5427;
    wire N__5424;
    wire N__5421;
    wire N__5418;
    wire N__5415;
    wire N__5412;
    wire N__5409;
    wire N__5406;
    wire N__5405;
    wire N__5404;
    wire N__5401;
    wire N__5400;
    wire N__5397;
    wire N__5394;
    wire N__5391;
    wire N__5388;
    wire N__5383;
    wire N__5380;
    wire N__5377;
    wire N__5374;
    wire N__5369;
    wire N__5364;
    wire N__5363;
    wire N__5358;
    wire N__5357;
    wire N__5356;
    wire N__5355;
    wire N__5352;
    wire N__5347;
    wire N__5344;
    wire N__5337;
    wire N__5336;
    wire N__5335;
    wire N__5332;
    wire N__5329;
    wire N__5328;
    wire N__5327;
    wire N__5324;
    wire N__5323;
    wire N__5322;
    wire N__5321;
    wire N__5320;
    wire N__5319;
    wire N__5316;
    wire N__5315;
    wire N__5312;
    wire N__5307;
    wire N__5304;
    wire N__5303;
    wire N__5302;
    wire N__5301;
    wire N__5298;
    wire N__5297;
    wire N__5296;
    wire N__5295;
    wire N__5294;
    wire N__5291;
    wire N__5284;
    wire N__5281;
    wire N__5278;
    wire N__5271;
    wire N__5260;
    wire N__5257;
    wire N__5252;
    wire N__5235;
    wire N__5234;
    wire N__5231;
    wire N__5228;
    wire N__5227;
    wire N__5226;
    wire N__5225;
    wire N__5224;
    wire N__5223;
    wire N__5222;
    wire N__5217;
    wire N__5214;
    wire N__5211;
    wire N__5210;
    wire N__5209;
    wire N__5208;
    wire N__5207;
    wire N__5206;
    wire N__5203;
    wire N__5202;
    wire N__5201;
    wire N__5200;
    wire N__5197;
    wire N__5194;
    wire N__5191;
    wire N__5186;
    wire N__5183;
    wire N__5170;
    wire N__5161;
    wire N__5148;
    wire N__5147;
    wire N__5146;
    wire N__5145;
    wire N__5144;
    wire N__5143;
    wire N__5142;
    wire N__5141;
    wire N__5134;
    wire N__5133;
    wire N__5132;
    wire N__5131;
    wire N__5130;
    wire N__5127;
    wire N__5122;
    wire N__5119;
    wire N__5118;
    wire N__5115;
    wire N__5112;
    wire N__5111;
    wire N__5108;
    wire N__5107;
    wire N__5106;
    wire N__5103;
    wire N__5102;
    wire N__5101;
    wire N__5100;
    wire N__5097;
    wire N__5094;
    wire N__5089;
    wire N__5086;
    wire N__5081;
    wire N__5078;
    wire N__5067;
    wire N__5064;
    wire N__5059;
    wire N__5040;
    wire N__5039;
    wire N__5038;
    wire N__5037;
    wire N__5034;
    wire N__5029;
    wire N__5026;
    wire N__5025;
    wire N__5024;
    wire N__5023;
    wire N__5022;
    wire N__5021;
    wire N__5020;
    wire N__5019;
    wire N__5018;
    wire N__5013;
    wire N__5010;
    wire N__5005;
    wire N__4992;
    wire N__4991;
    wire N__4990;
    wire N__4989;
    wire N__4988;
    wire N__4979;
    wire N__4970;
    wire N__4965;
    wire N__4964;
    wire N__4963;
    wire N__4960;
    wire N__4959;
    wire N__4956;
    wire N__4955;
    wire N__4952;
    wire N__4949;
    wire N__4946;
    wire N__4941;
    wire N__4938;
    wire N__4931;
    wire N__4926;
    wire N__4923;
    wire N__4920;
    wire N__4917;
    wire N__4916;
    wire N__4915;
    wire N__4912;
    wire N__4909;
    wire N__4906;
    wire N__4903;
    wire N__4902;
    wire N__4901;
    wire N__4898;
    wire N__4895;
    wire N__4892;
    wire N__4887;
    wire N__4878;
    wire N__4875;
    wire N__4872;
    wire N__4871;
    wire N__4868;
    wire N__4865;
    wire N__4862;
    wire N__4859;
    wire N__4854;
    wire N__4851;
    wire N__4848;
    wire N__4845;
    wire N__4842;
    wire N__4839;
    wire N__4836;
    wire N__4833;
    wire N__4830;
    wire N__4829;
    wire N__4826;
    wire N__4823;
    wire N__4818;
    wire N__4815;
    wire N__4812;
    wire N__4809;
    wire N__4808;
    wire N__4807;
    wire N__4806;
    wire N__4805;
    wire N__4802;
    wire N__4797;
    wire N__4794;
    wire N__4791;
    wire N__4790;
    wire N__4789;
    wire N__4782;
    wire N__4781;
    wire N__4774;
    wire N__4771;
    wire N__4768;
    wire N__4761;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4746;
    wire N__4743;
    wire N__4740;
    wire N__4737;
    wire N__4734;
    wire N__4731;
    wire N__4728;
    wire N__4725;
    wire N__4724;
    wire N__4719;
    wire N__4716;
    wire N__4713;
    wire N__4710;
    wire N__4707;
    wire N__4704;
    wire N__4701;
    wire N__4698;
    wire N__4697;
    wire N__4694;
    wire N__4691;
    wire N__4686;
    wire N__4685;
    wire N__4680;
    wire N__4677;
    wire N__4674;
    wire N__4671;
    wire N__4668;
    wire N__4665;
    wire N__4662;
    wire N__4659;
    wire N__4656;
    wire N__4653;
    wire N__4650;
    wire N__4647;
    wire N__4644;
    wire N__4643;
    wire N__4638;
    wire N__4635;
    wire N__4632;
    wire N__4629;
    wire N__4626;
    wire N__4625;
    wire N__4624;
    wire N__4623;
    wire N__4622;
    wire N__4621;
    wire N__4620;
    wire N__4617;
    wire N__4614;
    wire N__4607;
    wire N__4606;
    wire N__4605;
    wire N__4604;
    wire N__4599;
    wire N__4594;
    wire N__4591;
    wire N__4588;
    wire N__4583;
    wire N__4582;
    wire N__4581;
    wire N__4580;
    wire N__4579;
    wire N__4578;
    wire N__4575;
    wire N__4570;
    wire N__4567;
    wire N__4564;
    wire N__4557;
    wire N__4552;
    wire N__4539;
    wire N__4538;
    wire N__4535;
    wire N__4532;
    wire N__4527;
    wire N__4524;
    wire N__4521;
    wire N__4520;
    wire N__4517;
    wire N__4514;
    wire N__4509;
    wire N__4508;
    wire N__4503;
    wire N__4500;
    wire N__4497;
    wire N__4494;
    wire N__4491;
    wire N__4490;
    wire N__4487;
    wire N__4484;
    wire N__4481;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4469;
    wire N__4466;
    wire N__4461;
    wire N__4460;
    wire N__4459;
    wire N__4456;
    wire N__4455;
    wire N__4454;
    wire N__4453;
    wire N__4450;
    wire N__4447;
    wire N__4442;
    wire N__4439;
    wire N__4438;
    wire N__4435;
    wire N__4432;
    wire N__4429;
    wire N__4426;
    wire N__4423;
    wire N__4420;
    wire N__4419;
    wire N__4418;
    wire N__4415;
    wire N__4410;
    wire N__4405;
    wire N__4398;
    wire N__4389;
    wire N__4388;
    wire N__4387;
    wire N__4386;
    wire N__4385;
    wire N__4384;
    wire N__4377;
    wire N__4372;
    wire N__4369;
    wire N__4366;
    wire N__4363;
    wire N__4362;
    wire N__4361;
    wire N__4360;
    wire N__4359;
    wire N__4356;
    wire N__4353;
    wire N__4350;
    wire N__4341;
    wire N__4332;
    wire N__4331;
    wire N__4328;
    wire N__4327;
    wire N__4324;
    wire N__4323;
    wire N__4322;
    wire N__4321;
    wire N__4318;
    wire N__4315;
    wire N__4312;
    wire N__4307;
    wire N__4304;
    wire N__4301;
    wire N__4298;
    wire N__4295;
    wire N__4292;
    wire N__4281;
    wire N__4278;
    wire N__4275;
    wire N__4272;
    wire N__4269;
    wire N__4266;
    wire N__4263;
    wire N__4260;
    wire N__4257;
    wire N__4254;
    wire N__4251;
    wire N__4248;
    wire N__4245;
    wire N__4242;
    wire N__4239;
    wire N__4238;
    wire N__4235;
    wire N__4232;
    wire N__4231;
    wire N__4230;
    wire N__4227;
    wire N__4224;
    wire N__4223;
    wire N__4220;
    wire N__4217;
    wire N__4214;
    wire N__4211;
    wire N__4204;
    wire N__4197;
    wire N__4194;
    wire N__4191;
    wire N__4188;
    wire N__4187;
    wire N__4184;
    wire N__4183;
    wire N__4182;
    wire N__4179;
    wire N__4178;
    wire N__4177;
    wire N__4174;
    wire N__4171;
    wire N__4164;
    wire N__4161;
    wire N__4160;
    wire N__4157;
    wire N__4154;
    wire N__4151;
    wire N__4146;
    wire N__4137;
    wire N__4134;
    wire N__4133;
    wire N__4130;
    wire N__4129;
    wire N__4126;
    wire N__4123;
    wire N__4120;
    wire N__4117;
    wire N__4114;
    wire N__4107;
    wire N__4106;
    wire N__4103;
    wire N__4100;
    wire N__4095;
    wire N__4092;
    wire N__4089;
    wire N__4086;
    wire N__4085;
    wire N__4080;
    wire N__4077;
    wire N__4074;
    wire N__4071;
    wire N__4068;
    wire N__4065;
    wire N__4062;
    wire N__4059;
    wire N__4056;
    wire N__4053;
    wire N__4050;
    wire N__4047;
    wire N__4044;
    wire N__4041;
    wire N__4038;
    wire N__4037;
    wire N__4036;
    wire N__4033;
    wire N__4028;
    wire N__4025;
    wire N__4020;
    wire N__4017;
    wire N__4014;
    wire N__4011;
    wire N__4008;
    wire N__4005;
    wire N__4002;
    wire N__3999;
    wire N__3996;
    wire N__3993;
    wire N__3990;
    wire N__3987;
    wire N__3984;
    wire N__3983;
    wire N__3982;
    wire N__3979;
    wire N__3976;
    wire N__3973;
    wire N__3970;
    wire N__3963;
    wire N__3960;
    wire N__3957;
    wire N__3954;
    wire N__3951;
    wire N__3948;
    wire N__3945;
    wire N__3942;
    wire N__3939;
    wire N__3936;
    wire N__3933;
    wire N__3930;
    wire N__3929;
    wire N__3926;
    wire N__3923;
    wire N__3918;
    wire N__3915;
    wire N__3912;
    wire N__3909;
    wire N__3906;
    wire N__3903;
    wire N__3900;
    wire N__3897;
    wire N__3894;
    wire N__3891;
    wire N__3888;
    wire N__3887;
    wire N__3886;
    wire N__3885;
    wire N__3884;
    wire N__3883;
    wire N__3882;
    wire N__3881;
    wire N__3880;
    wire N__3879;
    wire N__3864;
    wire N__3861;
    wire N__3858;
    wire N__3855;
    wire N__3846;
    wire N__3843;
    wire N__3842;
    wire N__3839;
    wire N__3836;
    wire N__3833;
    wire N__3830;
    wire N__3825;
    wire N__3822;
    wire N__3819;
    wire N__3816;
    wire N__3813;
    wire N__3810;
    wire N__3807;
    wire N__3804;
    wire N__3801;
    wire N__3798;
    wire N__3795;
    wire N__3792;
    wire N__3789;
    wire N__3786;
    wire N__3783;
    wire N__3780;
    wire N__3777;
    wire N__3774;
    wire N__3773;
    wire N__3772;
    wire N__3771;
    wire N__3770;
    wire N__3769;
    wire N__3768;
    wire N__3765;
    wire N__3754;
    wire N__3751;
    wire N__3746;
    wire N__3741;
    wire N__3740;
    wire N__3739;
    wire N__3738;
    wire N__3737;
    wire N__3736;
    wire N__3733;
    wire N__3722;
    wire N__3721;
    wire N__3716;
    wire N__3713;
    wire N__3708;
    wire N__3707;
    wire N__3706;
    wire N__3705;
    wire N__3702;
    wire N__3699;
    wire N__3696;
    wire N__3695;
    wire N__3692;
    wire N__3691;
    wire N__3688;
    wire N__3677;
    wire N__3676;
    wire N__3671;
    wire N__3668;
    wire N__3663;
    wire N__3662;
    wire N__3661;
    wire N__3660;
    wire N__3659;
    wire N__3656;
    wire N__3655;
    wire N__3652;
    wire N__3651;
    wire N__3648;
    wire N__3637;
    wire N__3634;
    wire N__3629;
    wire N__3626;
    wire N__3621;
    wire N__3618;
    wire N__3615;
    wire N__3612;
    wire N__3609;
    wire N__3606;
    wire N__3603;
    wire N__3600;
    wire N__3597;
    wire N__3594;
    wire N__3591;
    wire N__3588;
    wire N__3585;
    wire N__3582;
    wire N__3579;
    wire N__3576;
    wire N__3573;
    wire N__3570;
    wire N__3567;
    wire N__3566;
    wire N__3565;
    wire N__3562;
    wire N__3559;
    wire N__3556;
    wire N__3553;
    wire N__3546;
    wire N__3543;
    wire N__3542;
    wire N__3541;
    wire N__3538;
    wire N__3535;
    wire N__3532;
    wire N__3525;
    wire N__3522;
    wire N__3521;
    wire N__3518;
    wire N__3517;
    wire N__3514;
    wire N__3511;
    wire N__3508;
    wire N__3501;
    wire N__3498;
    wire N__3495;
    wire N__3494;
    wire N__3493;
    wire N__3490;
    wire N__3487;
    wire N__3484;
    wire N__3477;
    wire N__3474;
    wire N__3473;
    wire N__3472;
    wire N__3471;
    wire N__3468;
    wire N__3465;
    wire N__3462;
    wire N__3459;
    wire N__3456;
    wire N__3447;
    wire N__3446;
    wire N__3445;
    wire N__3444;
    wire N__3435;
    wire N__3432;
    wire N__3429;
    wire N__3426;
    wire N__3423;
    wire N__3420;
    wire N__3417;
    wire N__3414;
    wire N__3411;
    wire N__3410;
    wire N__3409;
    wire N__3406;
    wire N__3401;
    wire N__3396;
    wire N__3393;
    wire N__3392;
    wire N__3391;
    wire N__3388;
    wire N__3385;
    wire N__3380;
    wire N__3375;
    wire N__3372;
    wire N__3369;
    wire N__3368;
    wire N__3367;
    wire N__3364;
    wire N__3359;
    wire N__3354;
    wire N__3351;
    wire N__3350;
    wire N__3349;
    wire N__3346;
    wire N__3343;
    wire N__3340;
    wire N__3337;
    wire N__3330;
    wire N__3327;
    wire N__3324;
    wire N__3323;
    wire N__3322;
    wire N__3319;
    wire N__3316;
    wire N__3313;
    wire N__3306;
    wire N__3303;
    wire N__3302;
    wire N__3301;
    wire N__3298;
    wire N__3295;
    wire N__3292;
    wire N__3285;
    wire N__3282;
    wire N__3281;
    wire N__3278;
    wire N__3277;
    wire N__3274;
    wire N__3269;
    wire N__3264;
    wire N__3261;
    wire N__3260;
    wire N__3259;
    wire N__3256;
    wire N__3251;
    wire N__3246;
    wire N__3243;
    wire N__3240;
    wire N__3237;
    wire N__3234;
    wire N__3231;
    wire N__3228;
    wire N__3225;
    wire N__3222;
    wire N__3221;
    wire N__3220;
    wire N__3217;
    wire N__3212;
    wire N__3207;
    wire N__3206;
    wire N__3203;
    wire N__3200;
    wire N__3195;
    wire N__3192;
    wire N__3191;
    wire N__3188;
    wire N__3185;
    wire N__3182;
    wire N__3177;
    wire N__3174;
    wire N__3173;
    wire N__3172;
    wire N__3169;
    wire N__3166;
    wire N__3163;
    wire N__3158;
    wire N__3153;
    wire N__3150;
    wire N__3147;
    wire N__3146;
    wire N__3145;
    wire N__3142;
    wire N__3139;
    wire N__3136;
    wire N__3129;
    wire N__3126;
    wire N__3123;
    wire N__3120;
    wire N__3117;
    wire N__3114;
    wire N__3111;
    wire N__3108;
    wire N__3105;
    wire N__3102;
    wire N__3099;
    wire N__3096;
    wire N__3093;
    wire N__3090;
    wire N__3087;
    wire N__3084;
    wire N__3081;
    wire N__3078;
    wire N__3075;
    wire N__3072;
    wire N__3069;
    wire N__3066;
    wire N__3063;
    wire N__3060;
    wire N__3057;
    wire N__3054;
    wire N__3053;
    wire N__3050;
    wire N__3047;
    wire N__3044;
    wire N__3041;
    wire N__3038;
    wire N__3033;
    wire N__3030;
    wire N__3027;
    wire N__3024;
    wire N__3021;
    wire N__3018;
    wire N__3015;
    wire N__3014;
    wire N__3013;
    wire N__3012;
    wire N__3009;
    wire N__3002;
    wire N__2997;
    wire N__2994;
    wire N__2991;
    wire N__2988;
    wire N__2985;
    wire N__2982;
    wire GNDG0;
    wire VCCG0;
    wire \Instance1.un1_r_Count_10lt11_0_cascade_ ;
    wire \Instance1.un1_r_Count_10lto11_1 ;
    wire \Instance1.un1_r_Count_10lt17_cascade_ ;
    wire \Instance1.r_Count12_i ;
    wire \Instance1.un1_r_Count_10lto17_1 ;
    wire r_SwitchZ0Z_1;
    wire \Instance1.r_Count13_8_0 ;
    wire \Instance1.r_Count13_4_cascade_ ;
    wire \Instance1.r_Count13_7 ;
    wire \Instance1.r_Count13_10 ;
    wire i_Switch_1_c;
    wire \Instance1.r_Count13_12 ;
    wire \Instance1.r_Count13_13_cascade_ ;
    wire w_Switch_1;
    wire sevsegl_RNO_0Z0Z_2_cascade_;
    wire sevsegl_RNO_1Z0Z_2;
    wire r_HexEncode_i_0_6;
    wire r_HexEncode_i_1;
    wire r_HexEncode_i_0_5;
    wire SUM_2;
    wire SUM_2_cascade_;
    wire r_HexEncode_i_0_0;
    wire r_HexEncode_i_0_1;
    wire r_HexEncode_i_6;
    wire \Instance1.r_CountZ0Z_1 ;
    wire bfn_2_9_0_;
    wire \Instance1.r_CountZ0Z_2 ;
    wire \Instance1.r_Count_2_cry_1 ;
    wire \Instance1.r_CountZ0Z_3 ;
    wire \Instance1.r_Count_2_cry_2 ;
    wire \Instance1.r_CountZ0Z_4 ;
    wire \Instance1.r_Count_2_cry_3 ;
    wire \Instance1.r_CountZ0Z_5 ;
    wire \Instance1.r_Count_2_cry_4 ;
    wire \Instance1.r_CountZ0Z_6 ;
    wire \Instance1.r_Count_2_cry_5 ;
    wire \Instance1.r_CountZ0Z_7 ;
    wire \Instance1.r_Count_2_cry_6 ;
    wire \Instance1.r_CountZ0Z_8 ;
    wire \Instance1.r_Count_2_cry_7 ;
    wire \Instance1.r_Count_2_cry_8 ;
    wire \Instance1.r_CountZ0Z_9 ;
    wire bfn_2_10_0_;
    wire \Instance1.r_CountZ0Z_10 ;
    wire \Instance1.r_Count_2_cry_9 ;
    wire \Instance1.r_CountZ0Z_11 ;
    wire \Instance1.r_Count_2_cry_10 ;
    wire \Instance1.r_CountZ0Z_12 ;
    wire \Instance1.r_Count_2_cry_11 ;
    wire \Instance1.r_CountZ0Z_13 ;
    wire \Instance1.r_Count_2_cry_12 ;
    wire \Instance1.r_CountZ0Z_14 ;
    wire \Instance1.r_Count_2_cry_13 ;
    wire \Instance1.r_CountZ0Z_15 ;
    wire \Instance1.r_Count_2_cry_14 ;
    wire \Instance1.r_CountZ0Z_16 ;
    wire \Instance1.r_Count_2_cry_15 ;
    wire \Instance1.r_Count_2_cry_16 ;
    wire bfn_2_11_0_;
    wire \Instance1.r_CountZ0Z_17 ;
    wire \Instance1.r_CountZ0Z_0 ;
    wire \Instance1.r_Count12_i_g ;
    wire left_1;
    wire right_1;
    wire sevsegl_RNO_1Z0Z_3;
    wire sevsegr_RNO_1Z0Z_1;
    wire sevsegr_RNO_1Z0Z_2;
    wire sevsegr_RNO_0Z0Z_3;
    wire sevsegl_RNO_1Z0Z_1;
    wire sevsegr_7_ns_1_0;
    wire sevsegl_7_ns_1_0;
    wire r_Switch_2_RNIK7AZ0Z11;
    wire un1_click17_0;
    wire r_HexEncode_i_4;
    wire r_HexEncode_i_0;
    wire r_HexEncode_i_2;
    wire r_HexEncode_i_3;
    wire sevsegrZ0Z_0;
    wire sevsegrZ0Z_2;
    wire sevsegrZ0Z_1;
    wire sevsegrZ0Z_3;
    wire r_HexEncode_i_5;
    wire SUM_3_cascade_;
    wire r_Count11;
    wire r_Count11_cascade_;
    wire \alogicunit.N_95_1_cascade_ ;
    wire right_0;
    wire right_3;
    wire SUM_3;
    wire sevsegr_RNO_1Z0Z_3;
    wire right_2;
    wire bfn_4_12_0_;
    wire \alogicunit.un1_a_1_cry_1_THRU_CO ;
    wire \alogicunit.un1_a_1_cry_1 ;
    wire \alogicunit.un1_a_1_cry_2_THRU_CO ;
    wire \alogicunit.un1_a_1_cry_2 ;
    wire \alogicunit.un1_a_1_cry_3 ;
    wire \alogicunit.result_RNO_0Z0Z_5 ;
    wire \alogicunit.un1_a_1_cry_4 ;
    wire \alogicunit.un1_a_1_cry_5 ;
    wire \alogicunit.N_95_1 ;
    wire \alogicunit.un1_a_1_cry_6 ;
    wire left_3;
    wire \alogicunit.m26_l_fxZ0Z_0 ;
    wire un1_click13_1_sn_cascade_;
    wire sevsegr_RNO_0Z0Z_2;
    wire sevsegr_RNO_0Z0Z_1;
    wire r_SwitchZ0Z_3;
    wire \alogicunit.m26_l_fxZ0 ;
    wire sevsegl_RNO_0Z0Z_1;
    wire r_CountZ0Z_3;
    wire sevsegl_RNO_0Z0Z_3;
    wire \alogicunit.result24 ;
    wire \alogicunit.result24_cascade_ ;
    wire \alogicunit.un1_a_1_axb_3 ;
    wire \alogicunit.N_51 ;
    wire cu1_track_ns_3;
    wire N_28;
    wire \alogicunit.N_41 ;
    wire \alogicunit.N_41_cascade_ ;
    wire track_RNI9MAL_0_1;
    wire r_CountZ0Z_1;
    wire r_CountZ0Z_0;
    wire r_CountZ0Z_2;
    wire \Instance2.r_Count13_8_0_cascade_ ;
    wire \Instance2.un1_r_Count_10lt11_0_cascade_ ;
    wire \Instance2.r_Count13_12 ;
    wire \Instance2.r_Count13_13_cascade_ ;
    wire \Instance2.un1_r_Count_10lto11_1 ;
    wire \Instance2.r_Count13_10 ;
    wire \Instance2.r_Count13_7 ;
    wire \alogicunit.N_90 ;
    wire \Instance2.r_Count13_4 ;
    wire click13;
    wire \alogicunit.N_49 ;
    wire r_SwitchZ0Z_2;
    wire r_SwitchZ0Z_4;
    wire \Instance2.click14_sn_cascade_ ;
    wire un1_click13_1_sn;
    wire Instance2_un1_click13_3_1;
    wire \alogicunit.result_RNO_0Z0Z_4 ;
    wire left_0;
    wire \alogicunit.N_50 ;
    wire \alogicunit.result_RNO_0Z0Z_6 ;
    wire left_2;
    wire \alogicunit.un1_a_1_cry_1_c_invZ0 ;
    wire \alogicunit.N_102 ;
    wire r_HexEncode_i_0_4;
    wire \alogicunit.N_35 ;
    wire \alogicunit.result24_iZ0 ;
    wire current_state_0;
    wire current_state_1;
    wire current_state_2;
    wire current_state_3;
    wire clickZ0Z1;
    wire \Instance2.un1_r_Count_10lto17_1 ;
    wire w_Switch_2;
    wire i_Switch_2_c;
    wire \Instance2.un1_r_Count_10lt17 ;
    wire \Instance2.r_Count12_i ;
    wire bfn_6_7_0_;
    wire \Instance4.r_Count_2_cry_1 ;
    wire \Instance4.r_Count_2_cry_2 ;
    wire \Instance4.r_Count_2_cry_3 ;
    wire \Instance4.r_Count_2_cry_4 ;
    wire \Instance4.r_Count_2_cry_5 ;
    wire \Instance4.r_Count_2_cry_6 ;
    wire \Instance4.r_Count_2_cry_7 ;
    wire \Instance4.r_Count_2_cry_8 ;
    wire bfn_6_8_0_;
    wire \Instance4.r_Count_2_cry_9 ;
    wire \Instance4.r_Count_2_cry_10 ;
    wire \Instance4.r_Count_2_cry_11 ;
    wire \Instance4.r_Count_2_cry_12 ;
    wire \Instance4.r_Count_2_cry_13 ;
    wire \Instance4.r_Count_2_cry_14 ;
    wire \Instance4.r_Count_2_cry_15 ;
    wire \Instance4.r_Count_2_cry_16 ;
    wire bfn_6_9_0_;
    wire \Instance4.r_Count12_i_g ;
    wire bfn_6_10_0_;
    wire \Instance2.r_Count_0_2 ;
    wire \Instance2.r_Count_2_cry_1 ;
    wire \Instance2.r_Count_0_3 ;
    wire \Instance2.r_Count_2_cry_2 ;
    wire \Instance2.r_CountZ0Z_4 ;
    wire \Instance2.r_Count_2_cry_3 ;
    wire \Instance2.r_CountZ0Z_5 ;
    wire \Instance2.r_Count_2_cry_4 ;
    wire \Instance2.r_CountZ0Z_6 ;
    wire \Instance2.r_Count_2_cry_5 ;
    wire \Instance2.r_CountZ0Z_7 ;
    wire \Instance2.r_Count_2_cry_6 ;
    wire \Instance2.r_CountZ0Z_8 ;
    wire \Instance2.r_Count_2_cry_7 ;
    wire \Instance2.r_Count_2_cry_8 ;
    wire \Instance2.r_CountZ0Z_9 ;
    wire bfn_6_11_0_;
    wire \Instance2.r_CountZ0Z_10 ;
    wire \Instance2.r_Count_2_cry_9 ;
    wire \Instance2.r_CountZ0Z_11 ;
    wire \Instance2.r_Count_2_cry_10 ;
    wire \Instance2.r_CountZ0Z_12 ;
    wire \Instance2.r_Count_2_cry_11 ;
    wire \Instance2.r_CountZ0Z_13 ;
    wire \Instance2.r_Count_2_cry_12 ;
    wire \Instance2.r_CountZ0Z_14 ;
    wire \Instance2.r_Count_2_cry_13 ;
    wire \Instance2.r_CountZ0Z_15 ;
    wire \Instance2.r_Count_2_cry_14 ;
    wire \Instance2.r_CountZ0Z_16 ;
    wire \Instance2.r_Count_2_cry_15 ;
    wire \Instance2.r_Count_2_cry_16 ;
    wire bfn_6_12_0_;
    wire \Instance2.r_CountZ0Z_17 ;
    wire \Instance2.r_Count_0_0 ;
    wire \Instance2.r_Count_0_1 ;
    wire \Instance2.r_Count12_i_g ;
    wire CONSTANT_ONE_NET;
    wire r_HexEncode_i_0_3;
    wire sevseglZ0Z_2;
    wire sevseglZ0Z_1;
    wire sevseglZ0Z_3;
    wire sevseglZ0Z_0;
    wire r_HexEncode_i_0_2;
    wire \Instance4.r_CountZ0Z_1 ;
    wire \Instance4.r_CountZ0Z_2 ;
    wire \Instance4.r_CountZ0Z_3 ;
    wire \Instance4.r_CountZ0Z_4 ;
    wire \Instance4.r_CountZ0Z_7 ;
    wire \Instance4.r_CountZ0Z_0 ;
    wire \Instance4.r_Count13_8_0_cascade_ ;
    wire \Instance4.r_CountZ0Z_5 ;
    wire \Instance4.r_Count13_7 ;
    wire \Instance4.r_Count13_13_cascade_ ;
    wire \Instance4.r_Count13_12 ;
    wire \Instance4.r_CountZ0Z_14 ;
    wire \Instance4.r_CountZ0Z_17 ;
    wire \Instance4.r_Count13_4 ;
    wire \Instance4.r_CountZ0Z_11 ;
    wire \Instance4.r_CountZ0Z_10 ;
    wire \Instance4.r_CountZ0Z_9 ;
    wire \Instance4.r_CountZ0Z_13 ;
    wire \Instance4.r_CountZ0Z_12 ;
    wire \Instance4.un1_r_Count_10lto11_1_cascade_ ;
    wire \Instance4.un1_r_Count_10lt11_0 ;
    wire i_Switch_4_c;
    wire w_Switch_4;
    wire \Instance4.un1_r_Count_10lt17_cascade_ ;
    wire \Instance4.un1_r_Count_10lto17_1 ;
    wire \Instance4.r_Count12_i ;
    wire \Instance4.r_CountZ0Z_8 ;
    wire \Instance4.r_CountZ0Z_15 ;
    wire \Instance4.r_CountZ0Z_16 ;
    wire \Instance4.r_CountZ0Z_6 ;
    wire \Instance4.r_Count13_10 ;
    wire w_Switch_3;
    wire i_Switch_3_c;
    wire \Instance3.un1_r_Count_10lt17_cascade_ ;
    wire \Instance3.r_Count12_i ;
    wire \Instance3.r_Count13_8_0_cascade_ ;
    wire \Instance3.r_Count13_12 ;
    wire \Instance3.un1_r_Count_10lt11_0 ;
    wire \Instance3.un1_r_Count_10lto11_1 ;
    wire \Instance3.r_Count13_4 ;
    wire \Instance3.r_Count13_7_cascade_ ;
    wire \Instance3.r_Count13_13 ;
    wire \Instance3.r_Count13_10 ;
    wire \Instance3.un1_r_Count_10lto17_1 ;
    wire negative;
    wire o_LED_1_c;
    wire bfn_8_9_0_;
    wire \Instance3.r_CountZ0Z_2 ;
    wire \Instance3.r_Count_2_cry_1 ;
    wire \Instance3.r_CountZ0Z_3 ;
    wire \Instance3.r_Count_2_cry_2 ;
    wire \Instance3.r_CountZ0Z_4 ;
    wire \Instance3.r_Count_2_cry_3 ;
    wire \Instance3.r_CountZ0Z_5 ;
    wire \Instance3.r_Count_2_cry_4 ;
    wire \Instance3.r_CountZ0Z_6 ;
    wire \Instance3.r_Count_2_cry_5 ;
    wire \Instance3.r_CountZ0Z_7 ;
    wire \Instance3.r_Count_2_cry_6 ;
    wire \Instance3.r_CountZ0Z_8 ;
    wire \Instance3.r_Count_2_cry_7 ;
    wire \Instance3.r_Count_2_cry_8 ;
    wire \Instance3.r_CountZ0Z_9 ;
    wire bfn_8_10_0_;
    wire \Instance3.r_CountZ0Z_10 ;
    wire \Instance3.r_Count_2_cry_9 ;
    wire \Instance3.r_CountZ0Z_11 ;
    wire \Instance3.r_Count_2_cry_10 ;
    wire \Instance3.r_CountZ0Z_12 ;
    wire \Instance3.r_Count_2_cry_11 ;
    wire \Instance3.r_CountZ0Z_13 ;
    wire \Instance3.r_Count_2_cry_12 ;
    wire \Instance3.r_CountZ0Z_14 ;
    wire \Instance3.r_Count_2_cry_13 ;
    wire \Instance3.r_CountZ0Z_15 ;
    wire \Instance3.r_Count_2_cry_14 ;
    wire \Instance3.r_CountZ0Z_16 ;
    wire \Instance3.r_Count_2_cry_15 ;
    wire \Instance3.r_Count_2_cry_16 ;
    wire bfn_8_11_0_;
    wire \Instance3.r_CountZ0Z_17 ;
    wire \Instance3.r_CountZ0Z_0 ;
    wire \Instance3.r_CountZ0Z_1 ;
    wire _gnd_net_;
    wire i_Clk_c_g;
    wire \Instance3.r_Count12_i_g ;

    PRE_IO_GBUF i_Clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__7468),
            .GLOBALBUFFEROUTPUT(i_Clk_c_g));
    IO_PAD i_Clk_ibuf_gb_io_iopad (
            .OE(N__7470),
            .DIN(N__7469),
            .DOUT(N__7468),
            .PACKAGEPIN(i_Clk));
    defparam i_Clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam i_Clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO i_Clk_ibuf_gb_io_preio (
            .PADOEN(N__7470),
            .PADOUT(N__7469),
            .PADIN(N__7468),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_F_obuf_iopad (
            .OE(N__7459),
            .DIN(N__7458),
            .DOUT(N__7457),
            .PACKAGEPIN(o_Segment2_F));
    defparam o_Segment2_F_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_F_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_F_obuf_preio (
            .PADOEN(N__7459),
            .PADOUT(N__7458),
            .PADIN(N__7457),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3111),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_1_obuf_iopad (
            .OE(N__7450),
            .DIN(N__7449),
            .DOUT(N__7448),
            .PACKAGEPIN(o_LED_1));
    defparam o_LED_1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_1_obuf_preio (
            .PADOEN(N__7450),
            .PADOUT(N__7449),
            .PADIN(N__7448),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6759),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment1_G_obuf_iopad (
            .OE(N__7441),
            .DIN(N__7440),
            .DOUT(N__7439),
            .PACKAGEPIN(o_Segment1_G));
    defparam o_Segment1_G_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment1_G_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment1_G_obuf_preio (
            .PADOEN(N__7441),
            .PADOUT(N__7440),
            .PADIN(N__7439),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3240),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD i_Switch_4_ibuf_iopad (
            .OE(N__7432),
            .DIN(N__7431),
            .DOUT(N__7430),
            .PACKAGEPIN(i_Switch_4));
    defparam i_Switch_4_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam i_Switch_4_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO i_Switch_4_ibuf_preio (
            .PADOEN(N__7432),
            .PADOUT(N__7431),
            .PADIN(N__7430),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(i_Switch_4_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD i_Switch_1_ibuf_iopad (
            .OE(N__7423),
            .DIN(N__7422),
            .DOUT(N__7421),
            .PACKAGEPIN(i_Switch_1));
    defparam i_Switch_1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam i_Switch_1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO i_Switch_1_ibuf_preio (
            .PADOEN(N__7423),
            .PADOUT(N__7422),
            .PADIN(N__7421),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(i_Switch_1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment1_B_obuf_iopad (
            .OE(N__7414),
            .DIN(N__7413),
            .DOUT(N__7412),
            .PACKAGEPIN(o_Segment1_B));
    defparam o_Segment1_B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment1_B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment1_B_obuf_preio (
            .PADOEN(N__7414),
            .PADOUT(N__7413),
            .PADIN(N__7412),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3105),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD i_Switch_3_ibuf_iopad (
            .OE(N__7405),
            .DIN(N__7404),
            .DOUT(N__7403),
            .PACKAGEPIN(i_Switch_3));
    defparam i_Switch_3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam i_Switch_3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO i_Switch_3_ibuf_preio (
            .PADOEN(N__7405),
            .PADOUT(N__7404),
            .PADIN(N__7403),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(i_Switch_3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment1_E_obuf_iopad (
            .OE(N__7396),
            .DIN(N__7395),
            .DOUT(N__7394),
            .PACKAGEPIN(o_Segment1_E));
    defparam o_Segment1_E_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment1_E_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment1_E_obuf_preio (
            .PADOEN(N__7396),
            .PADOUT(N__7395),
            .PADIN(N__7394),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5892),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_2_obuf_iopad (
            .OE(N__7387),
            .DIN(N__7386),
            .DOUT(N__7385),
            .PACKAGEPIN(o_LED_2));
    defparam o_LED_2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_2_obuf_preio (
            .PADOEN(N__7387),
            .PADOUT(N__7386),
            .PADIN(N__7385),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6757),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_E_obuf_iopad (
            .OE(N__7378),
            .DIN(N__7377),
            .DOUT(N__7376),
            .PACKAGEPIN(o_Segment2_E));
    defparam o_Segment2_E_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_E_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_E_obuf_preio (
            .PADOEN(N__7378),
            .PADOUT(N__7377),
            .PADIN(N__7376),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3804),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_C_obuf_iopad (
            .OE(N__7369),
            .DIN(N__7368),
            .DOUT(N__7367),
            .PACKAGEPIN(o_Segment2_C));
    defparam o_Segment2_C_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_C_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_C_obuf_preio (
            .PADOEN(N__7369),
            .PADOUT(N__7368),
            .PADIN(N__7367),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3825),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_4_obuf_iopad (
            .OE(N__7360),
            .DIN(N__7359),
            .DOUT(N__7358),
            .PACKAGEPIN(o_LED_4));
    defparam o_LED_4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_4_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_4_obuf_preio (
            .PADOEN(N__7360),
            .PADOUT(N__7359),
            .PADIN(N__7358),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6747),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment1_A_obuf_iopad (
            .OE(N__7351),
            .DIN(N__7350),
            .DOUT(N__7349),
            .PACKAGEPIN(o_Segment1_A));
    defparam o_Segment1_A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment1_A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment1_A_obuf_preio (
            .PADOEN(N__7351),
            .PADOUT(N__7350),
            .PADIN(N__7349),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3117),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD i_Switch_2_ibuf_iopad (
            .OE(N__7342),
            .DIN(N__7341),
            .DOUT(N__7340),
            .PACKAGEPIN(i_Switch_2));
    defparam i_Switch_2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam i_Switch_2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO i_Switch_2_ibuf_preio (
            .PADOEN(N__7342),
            .PADOUT(N__7341),
            .PADIN(N__7340),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(i_Switch_2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_B_obuf_iopad (
            .OE(N__7333),
            .DIN(N__7332),
            .DOUT(N__7331),
            .PACKAGEPIN(o_Segment2_B));
    defparam o_Segment2_B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_B_obuf_preio (
            .PADOEN(N__7333),
            .PADOUT(N__7332),
            .PADIN(N__7331),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3621),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment1_C_obuf_iopad (
            .OE(N__7324),
            .DIN(N__7323),
            .DOUT(N__7322),
            .PACKAGEPIN(o_Segment1_C));
    defparam o_Segment1_C_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment1_C_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment1_C_obuf_preio (
            .PADOEN(N__7324),
            .PADOUT(N__7323),
            .PADIN(N__7322),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5415),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment1_D_obuf_iopad (
            .OE(N__7315),
            .DIN(N__7314),
            .DOUT(N__7313),
            .PACKAGEPIN(o_Segment1_D));
    defparam o_Segment1_D_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment1_D_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment1_D_obuf_preio (
            .PADOEN(N__7315),
            .PADOUT(N__7314),
            .PADIN(N__7313),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6087),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment1_F_obuf_iopad (
            .OE(N__7306),
            .DIN(N__7305),
            .DOUT(N__7304),
            .PACKAGEPIN(o_Segment1_F));
    defparam o_Segment1_F_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment1_F_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment1_F_obuf_preio (
            .PADOEN(N__7306),
            .PADOUT(N__7305),
            .PADIN(N__7304),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3234),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_3_obuf_iopad (
            .OE(N__7297),
            .DIN(N__7296),
            .DOUT(N__7295),
            .PACKAGEPIN(o_LED_3));
    defparam o_LED_3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_3_obuf_preio (
            .PADOEN(N__7297),
            .PADOUT(N__7296),
            .PADIN(N__7295),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6758),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_A_obuf_iopad (
            .OE(N__7288),
            .DIN(N__7287),
            .DOUT(N__7286),
            .PACKAGEPIN(o_Segment2_A));
    defparam o_Segment2_A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_A_obuf_preio (
            .PADOEN(N__7288),
            .PADOUT(N__7287),
            .PADIN(N__7286),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3228),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_G_obuf_iopad (
            .OE(N__7279),
            .DIN(N__7278),
            .DOUT(N__7277),
            .PACKAGEPIN(o_Segment2_G));
    defparam o_Segment2_G_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_G_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_G_obuf_preio (
            .PADOEN(N__7279),
            .PADOUT(N__7278),
            .PADIN(N__7277),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3819),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_D_obuf_iopad (
            .OE(N__7270),
            .DIN(N__7269),
            .DOUT(N__7268),
            .PACKAGEPIN(o_Segment2_D));
    defparam o_Segment2_D_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_D_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_D_obuf_preio (
            .PADOEN(N__7270),
            .PADOUT(N__7269),
            .PADIN(N__7268),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3792),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__1682 (
            .O(N__7251),
            .I(N__7246));
    InMux I__1681 (
            .O(N__7250),
            .I(N__7243));
    InMux I__1680 (
            .O(N__7249),
            .I(N__7238));
    InMux I__1679 (
            .O(N__7246),
            .I(N__7238));
    LocalMux I__1678 (
            .O(N__7243),
            .I(\Instance3.r_CountZ0Z_14 ));
    LocalMux I__1677 (
            .O(N__7238),
            .I(\Instance3.r_CountZ0Z_14 ));
    InMux I__1676 (
            .O(N__7233),
            .I(\Instance3.r_Count_2_cry_13 ));
    CascadeMux I__1675 (
            .O(N__7230),
            .I(N__7226));
    InMux I__1674 (
            .O(N__7229),
            .I(N__7222));
    InMux I__1673 (
            .O(N__7226),
            .I(N__7219));
    InMux I__1672 (
            .O(N__7225),
            .I(N__7216));
    LocalMux I__1671 (
            .O(N__7222),
            .I(\Instance3.r_CountZ0Z_15 ));
    LocalMux I__1670 (
            .O(N__7219),
            .I(\Instance3.r_CountZ0Z_15 ));
    LocalMux I__1669 (
            .O(N__7216),
            .I(\Instance3.r_CountZ0Z_15 ));
    InMux I__1668 (
            .O(N__7209),
            .I(\Instance3.r_Count_2_cry_14 ));
    InMux I__1667 (
            .O(N__7206),
            .I(N__7201));
    InMux I__1666 (
            .O(N__7205),
            .I(N__7198));
    InMux I__1665 (
            .O(N__7204),
            .I(N__7195));
    LocalMux I__1664 (
            .O(N__7201),
            .I(\Instance3.r_CountZ0Z_16 ));
    LocalMux I__1663 (
            .O(N__7198),
            .I(\Instance3.r_CountZ0Z_16 ));
    LocalMux I__1662 (
            .O(N__7195),
            .I(\Instance3.r_CountZ0Z_16 ));
    InMux I__1661 (
            .O(N__7188),
            .I(\Instance3.r_Count_2_cry_15 ));
    InMux I__1660 (
            .O(N__7185),
            .I(bfn_8_11_0_));
    InMux I__1659 (
            .O(N__7182),
            .I(N__7177));
    InMux I__1658 (
            .O(N__7181),
            .I(N__7172));
    InMux I__1657 (
            .O(N__7180),
            .I(N__7172));
    LocalMux I__1656 (
            .O(N__7177),
            .I(\Instance3.r_CountZ0Z_17 ));
    LocalMux I__1655 (
            .O(N__7172),
            .I(\Instance3.r_CountZ0Z_17 ));
    InMux I__1654 (
            .O(N__7167),
            .I(N__7164));
    LocalMux I__1653 (
            .O(N__7164),
            .I(N__7158));
    CascadeMux I__1652 (
            .O(N__7163),
            .I(N__7155));
    InMux I__1651 (
            .O(N__7162),
            .I(N__7150));
    InMux I__1650 (
            .O(N__7161),
            .I(N__7150));
    Span4Mux_v I__1649 (
            .O(N__7158),
            .I(N__7147));
    InMux I__1648 (
            .O(N__7155),
            .I(N__7144));
    LocalMux I__1647 (
            .O(N__7150),
            .I(\Instance3.r_CountZ0Z_0 ));
    Odrv4 I__1646 (
            .O(N__7147),
            .I(\Instance3.r_CountZ0Z_0 ));
    LocalMux I__1645 (
            .O(N__7144),
            .I(\Instance3.r_CountZ0Z_0 ));
    InMux I__1644 (
            .O(N__7137),
            .I(N__7132));
    InMux I__1643 (
            .O(N__7136),
            .I(N__7129));
    InMux I__1642 (
            .O(N__7135),
            .I(N__7126));
    LocalMux I__1641 (
            .O(N__7132),
            .I(N__7123));
    LocalMux I__1640 (
            .O(N__7129),
            .I(\Instance3.r_CountZ0Z_1 ));
    LocalMux I__1639 (
            .O(N__7126),
            .I(\Instance3.r_CountZ0Z_1 ));
    Odrv4 I__1638 (
            .O(N__7123),
            .I(\Instance3.r_CountZ0Z_1 ));
    ClkMux I__1637 (
            .O(N__7116),
            .I(N__7008));
    ClkMux I__1636 (
            .O(N__7115),
            .I(N__7008));
    ClkMux I__1635 (
            .O(N__7114),
            .I(N__7008));
    ClkMux I__1634 (
            .O(N__7113),
            .I(N__7008));
    ClkMux I__1633 (
            .O(N__7112),
            .I(N__7008));
    ClkMux I__1632 (
            .O(N__7111),
            .I(N__7008));
    ClkMux I__1631 (
            .O(N__7110),
            .I(N__7008));
    ClkMux I__1630 (
            .O(N__7109),
            .I(N__7008));
    ClkMux I__1629 (
            .O(N__7108),
            .I(N__7008));
    ClkMux I__1628 (
            .O(N__7107),
            .I(N__7008));
    ClkMux I__1627 (
            .O(N__7106),
            .I(N__7008));
    ClkMux I__1626 (
            .O(N__7105),
            .I(N__7008));
    ClkMux I__1625 (
            .O(N__7104),
            .I(N__7008));
    ClkMux I__1624 (
            .O(N__7103),
            .I(N__7008));
    ClkMux I__1623 (
            .O(N__7102),
            .I(N__7008));
    ClkMux I__1622 (
            .O(N__7101),
            .I(N__7008));
    ClkMux I__1621 (
            .O(N__7100),
            .I(N__7008));
    ClkMux I__1620 (
            .O(N__7099),
            .I(N__7008));
    ClkMux I__1619 (
            .O(N__7098),
            .I(N__7008));
    ClkMux I__1618 (
            .O(N__7097),
            .I(N__7008));
    ClkMux I__1617 (
            .O(N__7096),
            .I(N__7008));
    ClkMux I__1616 (
            .O(N__7095),
            .I(N__7008));
    ClkMux I__1615 (
            .O(N__7094),
            .I(N__7008));
    ClkMux I__1614 (
            .O(N__7093),
            .I(N__7008));
    ClkMux I__1613 (
            .O(N__7092),
            .I(N__7008));
    ClkMux I__1612 (
            .O(N__7091),
            .I(N__7008));
    ClkMux I__1611 (
            .O(N__7090),
            .I(N__7008));
    ClkMux I__1610 (
            .O(N__7089),
            .I(N__7008));
    ClkMux I__1609 (
            .O(N__7088),
            .I(N__7008));
    ClkMux I__1608 (
            .O(N__7087),
            .I(N__7008));
    ClkMux I__1607 (
            .O(N__7086),
            .I(N__7008));
    ClkMux I__1606 (
            .O(N__7085),
            .I(N__7008));
    ClkMux I__1605 (
            .O(N__7084),
            .I(N__7008));
    ClkMux I__1604 (
            .O(N__7083),
            .I(N__7008));
    ClkMux I__1603 (
            .O(N__7082),
            .I(N__7008));
    ClkMux I__1602 (
            .O(N__7081),
            .I(N__7008));
    GlobalMux I__1601 (
            .O(N__7008),
            .I(N__7005));
    gio2CtrlBuf I__1600 (
            .O(N__7005),
            .I(i_Clk_c_g));
    SRMux I__1599 (
            .O(N__7002),
            .I(N__6990));
    SRMux I__1598 (
            .O(N__7001),
            .I(N__6990));
    SRMux I__1597 (
            .O(N__7000),
            .I(N__6990));
    SRMux I__1596 (
            .O(N__6999),
            .I(N__6990));
    GlobalMux I__1595 (
            .O(N__6990),
            .I(N__6987));
    gio2CtrlBuf I__1594 (
            .O(N__6987),
            .I(\Instance3.r_Count12_i_g ));
    InMux I__1593 (
            .O(N__6984),
            .I(\Instance3.r_Count_2_cry_4 ));
    CascadeMux I__1592 (
            .O(N__6981),
            .I(N__6976));
    InMux I__1591 (
            .O(N__6980),
            .I(N__6973));
    InMux I__1590 (
            .O(N__6979),
            .I(N__6970));
    InMux I__1589 (
            .O(N__6976),
            .I(N__6967));
    LocalMux I__1588 (
            .O(N__6973),
            .I(\Instance3.r_CountZ0Z_6 ));
    LocalMux I__1587 (
            .O(N__6970),
            .I(\Instance3.r_CountZ0Z_6 ));
    LocalMux I__1586 (
            .O(N__6967),
            .I(\Instance3.r_CountZ0Z_6 ));
    InMux I__1585 (
            .O(N__6960),
            .I(\Instance3.r_Count_2_cry_5 ));
    InMux I__1584 (
            .O(N__6957),
            .I(N__6952));
    InMux I__1583 (
            .O(N__6956),
            .I(N__6947));
    InMux I__1582 (
            .O(N__6955),
            .I(N__6947));
    LocalMux I__1581 (
            .O(N__6952),
            .I(\Instance3.r_CountZ0Z_7 ));
    LocalMux I__1580 (
            .O(N__6947),
            .I(\Instance3.r_CountZ0Z_7 ));
    InMux I__1579 (
            .O(N__6942),
            .I(\Instance3.r_Count_2_cry_6 ));
    InMux I__1578 (
            .O(N__6939),
            .I(N__6934));
    InMux I__1577 (
            .O(N__6938),
            .I(N__6931));
    InMux I__1576 (
            .O(N__6937),
            .I(N__6928));
    LocalMux I__1575 (
            .O(N__6934),
            .I(\Instance3.r_CountZ0Z_8 ));
    LocalMux I__1574 (
            .O(N__6931),
            .I(\Instance3.r_CountZ0Z_8 ));
    LocalMux I__1573 (
            .O(N__6928),
            .I(\Instance3.r_CountZ0Z_8 ));
    InMux I__1572 (
            .O(N__6921),
            .I(\Instance3.r_Count_2_cry_7 ));
    InMux I__1571 (
            .O(N__6918),
            .I(N__6913));
    InMux I__1570 (
            .O(N__6917),
            .I(N__6910));
    InMux I__1569 (
            .O(N__6916),
            .I(N__6907));
    LocalMux I__1568 (
            .O(N__6913),
            .I(\Instance3.r_CountZ0Z_9 ));
    LocalMux I__1567 (
            .O(N__6910),
            .I(\Instance3.r_CountZ0Z_9 ));
    LocalMux I__1566 (
            .O(N__6907),
            .I(\Instance3.r_CountZ0Z_9 ));
    InMux I__1565 (
            .O(N__6900),
            .I(bfn_8_10_0_));
    CascadeMux I__1564 (
            .O(N__6897),
            .I(N__6894));
    InMux I__1563 (
            .O(N__6894),
            .I(N__6889));
    InMux I__1562 (
            .O(N__6893),
            .I(N__6886));
    InMux I__1561 (
            .O(N__6892),
            .I(N__6883));
    LocalMux I__1560 (
            .O(N__6889),
            .I(N__6880));
    LocalMux I__1559 (
            .O(N__6886),
            .I(\Instance3.r_CountZ0Z_10 ));
    LocalMux I__1558 (
            .O(N__6883),
            .I(\Instance3.r_CountZ0Z_10 ));
    Odrv4 I__1557 (
            .O(N__6880),
            .I(\Instance3.r_CountZ0Z_10 ));
    InMux I__1556 (
            .O(N__6873),
            .I(\Instance3.r_Count_2_cry_9 ));
    InMux I__1555 (
            .O(N__6870),
            .I(N__6865));
    InMux I__1554 (
            .O(N__6869),
            .I(N__6862));
    InMux I__1553 (
            .O(N__6868),
            .I(N__6859));
    LocalMux I__1552 (
            .O(N__6865),
            .I(N__6856));
    LocalMux I__1551 (
            .O(N__6862),
            .I(\Instance3.r_CountZ0Z_11 ));
    LocalMux I__1550 (
            .O(N__6859),
            .I(\Instance3.r_CountZ0Z_11 ));
    Odrv4 I__1549 (
            .O(N__6856),
            .I(\Instance3.r_CountZ0Z_11 ));
    InMux I__1548 (
            .O(N__6849),
            .I(\Instance3.r_Count_2_cry_10 ));
    CascadeMux I__1547 (
            .O(N__6846),
            .I(N__6843));
    InMux I__1546 (
            .O(N__6843),
            .I(N__6838));
    InMux I__1545 (
            .O(N__6842),
            .I(N__6835));
    InMux I__1544 (
            .O(N__6841),
            .I(N__6832));
    LocalMux I__1543 (
            .O(N__6838),
            .I(N__6829));
    LocalMux I__1542 (
            .O(N__6835),
            .I(\Instance3.r_CountZ0Z_12 ));
    LocalMux I__1541 (
            .O(N__6832),
            .I(\Instance3.r_CountZ0Z_12 ));
    Odrv4 I__1540 (
            .O(N__6829),
            .I(\Instance3.r_CountZ0Z_12 ));
    InMux I__1539 (
            .O(N__6822),
            .I(\Instance3.r_Count_2_cry_11 ));
    CascadeMux I__1538 (
            .O(N__6819),
            .I(N__6815));
    InMux I__1537 (
            .O(N__6818),
            .I(N__6811));
    InMux I__1536 (
            .O(N__6815),
            .I(N__6806));
    InMux I__1535 (
            .O(N__6814),
            .I(N__6806));
    LocalMux I__1534 (
            .O(N__6811),
            .I(\Instance3.r_CountZ0Z_13 ));
    LocalMux I__1533 (
            .O(N__6806),
            .I(\Instance3.r_CountZ0Z_13 ));
    InMux I__1532 (
            .O(N__6801),
            .I(\Instance3.r_Count_2_cry_12 ));
    CascadeMux I__1531 (
            .O(N__6798),
            .I(\Instance3.r_Count13_7_cascade_ ));
    InMux I__1530 (
            .O(N__6795),
            .I(N__6792));
    LocalMux I__1529 (
            .O(N__6792),
            .I(N__6789));
    Span4Mux_v I__1528 (
            .O(N__6789),
            .I(N__6786));
    Odrv4 I__1527 (
            .O(N__6786),
            .I(\Instance3.r_Count13_13 ));
    InMux I__1526 (
            .O(N__6783),
            .I(N__6780));
    LocalMux I__1525 (
            .O(N__6780),
            .I(\Instance3.r_Count13_10 ));
    InMux I__1524 (
            .O(N__6777),
            .I(N__6774));
    LocalMux I__1523 (
            .O(N__6774),
            .I(\Instance3.un1_r_Count_10lto17_1 ));
    InMux I__1522 (
            .O(N__6771),
            .I(N__6768));
    LocalMux I__1521 (
            .O(N__6768),
            .I(N__6765));
    Span4Mux_h I__1520 (
            .O(N__6765),
            .I(N__6762));
    Odrv4 I__1519 (
            .O(N__6762),
            .I(negative));
    IoInMux I__1518 (
            .O(N__6759),
            .I(N__6754));
    IoInMux I__1517 (
            .O(N__6758),
            .I(N__6751));
    IoInMux I__1516 (
            .O(N__6757),
            .I(N__6748));
    LocalMux I__1515 (
            .O(N__6754),
            .I(N__6744));
    LocalMux I__1514 (
            .O(N__6751),
            .I(N__6739));
    LocalMux I__1513 (
            .O(N__6748),
            .I(N__6739));
    IoInMux I__1512 (
            .O(N__6747),
            .I(N__6736));
    Span4Mux_s3_h I__1511 (
            .O(N__6744),
            .I(N__6733));
    Span4Mux_s3_h I__1510 (
            .O(N__6739),
            .I(N__6730));
    LocalMux I__1509 (
            .O(N__6736),
            .I(N__6727));
    Odrv4 I__1508 (
            .O(N__6733),
            .I(o_LED_1_c));
    Odrv4 I__1507 (
            .O(N__6730),
            .I(o_LED_1_c));
    Odrv12 I__1506 (
            .O(N__6727),
            .I(o_LED_1_c));
    InMux I__1505 (
            .O(N__6720),
            .I(N__6716));
    InMux I__1504 (
            .O(N__6719),
            .I(N__6713));
    LocalMux I__1503 (
            .O(N__6716),
            .I(\Instance3.r_CountZ0Z_2 ));
    LocalMux I__1502 (
            .O(N__6713),
            .I(\Instance3.r_CountZ0Z_2 ));
    InMux I__1501 (
            .O(N__6708),
            .I(\Instance3.r_Count_2_cry_1 ));
    CascadeMux I__1500 (
            .O(N__6705),
            .I(N__6701));
    InMux I__1499 (
            .O(N__6704),
            .I(N__6698));
    InMux I__1498 (
            .O(N__6701),
            .I(N__6695));
    LocalMux I__1497 (
            .O(N__6698),
            .I(\Instance3.r_CountZ0Z_3 ));
    LocalMux I__1496 (
            .O(N__6695),
            .I(\Instance3.r_CountZ0Z_3 ));
    InMux I__1495 (
            .O(N__6690),
            .I(\Instance3.r_Count_2_cry_2 ));
    InMux I__1494 (
            .O(N__6687),
            .I(N__6682));
    InMux I__1493 (
            .O(N__6686),
            .I(N__6677));
    InMux I__1492 (
            .O(N__6685),
            .I(N__6677));
    LocalMux I__1491 (
            .O(N__6682),
            .I(\Instance3.r_CountZ0Z_4 ));
    LocalMux I__1490 (
            .O(N__6677),
            .I(\Instance3.r_CountZ0Z_4 ));
    InMux I__1489 (
            .O(N__6672),
            .I(\Instance3.r_Count_2_cry_3 ));
    InMux I__1488 (
            .O(N__6669),
            .I(N__6664));
    InMux I__1487 (
            .O(N__6668),
            .I(N__6661));
    InMux I__1486 (
            .O(N__6667),
            .I(N__6658));
    LocalMux I__1485 (
            .O(N__6664),
            .I(N__6655));
    LocalMux I__1484 (
            .O(N__6661),
            .I(\Instance3.r_CountZ0Z_5 ));
    LocalMux I__1483 (
            .O(N__6658),
            .I(\Instance3.r_CountZ0Z_5 ));
    Odrv4 I__1482 (
            .O(N__6655),
            .I(\Instance3.r_CountZ0Z_5 ));
    InMux I__1481 (
            .O(N__6648),
            .I(N__6643));
    InMux I__1480 (
            .O(N__6647),
            .I(N__6640));
    InMux I__1479 (
            .O(N__6646),
            .I(N__6637));
    LocalMux I__1478 (
            .O(N__6643),
            .I(\Instance4.r_CountZ0Z_8 ));
    LocalMux I__1477 (
            .O(N__6640),
            .I(\Instance4.r_CountZ0Z_8 ));
    LocalMux I__1476 (
            .O(N__6637),
            .I(\Instance4.r_CountZ0Z_8 ));
    InMux I__1475 (
            .O(N__6630),
            .I(N__6625));
    InMux I__1474 (
            .O(N__6629),
            .I(N__6622));
    InMux I__1473 (
            .O(N__6628),
            .I(N__6619));
    LocalMux I__1472 (
            .O(N__6625),
            .I(\Instance4.r_CountZ0Z_15 ));
    LocalMux I__1471 (
            .O(N__6622),
            .I(\Instance4.r_CountZ0Z_15 ));
    LocalMux I__1470 (
            .O(N__6619),
            .I(\Instance4.r_CountZ0Z_15 ));
    CascadeMux I__1469 (
            .O(N__6612),
            .I(N__6608));
    InMux I__1468 (
            .O(N__6611),
            .I(N__6604));
    InMux I__1467 (
            .O(N__6608),
            .I(N__6599));
    InMux I__1466 (
            .O(N__6607),
            .I(N__6599));
    LocalMux I__1465 (
            .O(N__6604),
            .I(\Instance4.r_CountZ0Z_16 ));
    LocalMux I__1464 (
            .O(N__6599),
            .I(\Instance4.r_CountZ0Z_16 ));
    InMux I__1463 (
            .O(N__6594),
            .I(N__6589));
    InMux I__1462 (
            .O(N__6593),
            .I(N__6586));
    InMux I__1461 (
            .O(N__6592),
            .I(N__6583));
    LocalMux I__1460 (
            .O(N__6589),
            .I(\Instance4.r_CountZ0Z_6 ));
    LocalMux I__1459 (
            .O(N__6586),
            .I(\Instance4.r_CountZ0Z_6 ));
    LocalMux I__1458 (
            .O(N__6583),
            .I(\Instance4.r_CountZ0Z_6 ));
    CascadeMux I__1457 (
            .O(N__6576),
            .I(N__6573));
    InMux I__1456 (
            .O(N__6573),
            .I(N__6570));
    LocalMux I__1455 (
            .O(N__6570),
            .I(\Instance4.r_Count13_10 ));
    InMux I__1454 (
            .O(N__6567),
            .I(N__6564));
    LocalMux I__1453 (
            .O(N__6564),
            .I(N__6561));
    Span4Mux_v I__1452 (
            .O(N__6561),
            .I(N__6557));
    InMux I__1451 (
            .O(N__6560),
            .I(N__6552));
    Span4Mux_h I__1450 (
            .O(N__6557),
            .I(N__6549));
    InMux I__1449 (
            .O(N__6556),
            .I(N__6544));
    InMux I__1448 (
            .O(N__6555),
            .I(N__6544));
    LocalMux I__1447 (
            .O(N__6552),
            .I(w_Switch_3));
    Odrv4 I__1446 (
            .O(N__6549),
            .I(w_Switch_3));
    LocalMux I__1445 (
            .O(N__6544),
            .I(w_Switch_3));
    CascadeMux I__1444 (
            .O(N__6537),
            .I(N__6534));
    InMux I__1443 (
            .O(N__6534),
            .I(N__6531));
    LocalMux I__1442 (
            .O(N__6531),
            .I(N__6527));
    InMux I__1441 (
            .O(N__6530),
            .I(N__6524));
    Span4Mux_v I__1440 (
            .O(N__6527),
            .I(N__6521));
    LocalMux I__1439 (
            .O(N__6524),
            .I(N__6518));
    Span4Mux_h I__1438 (
            .O(N__6521),
            .I(N__6515));
    Span4Mux_v I__1437 (
            .O(N__6518),
            .I(N__6512));
    IoSpan4Mux I__1436 (
            .O(N__6515),
            .I(N__6509));
    Span4Mux_h I__1435 (
            .O(N__6512),
            .I(N__6506));
    Odrv4 I__1434 (
            .O(N__6509),
            .I(i_Switch_3_c));
    Odrv4 I__1433 (
            .O(N__6506),
            .I(i_Switch_3_c));
    CascadeMux I__1432 (
            .O(N__6501),
            .I(\Instance3.un1_r_Count_10lt17_cascade_ ));
    IoInMux I__1431 (
            .O(N__6498),
            .I(N__6495));
    LocalMux I__1430 (
            .O(N__6495),
            .I(N__6492));
    Odrv12 I__1429 (
            .O(N__6492),
            .I(\Instance3.r_Count12_i ));
    CascadeMux I__1428 (
            .O(N__6489),
            .I(\Instance3.r_Count13_8_0_cascade_ ));
    InMux I__1427 (
            .O(N__6486),
            .I(N__6483));
    LocalMux I__1426 (
            .O(N__6483),
            .I(N__6480));
    Span4Mux_h I__1425 (
            .O(N__6480),
            .I(N__6477));
    Odrv4 I__1424 (
            .O(N__6477),
            .I(\Instance3.r_Count13_12 ));
    InMux I__1423 (
            .O(N__6474),
            .I(N__6471));
    LocalMux I__1422 (
            .O(N__6471),
            .I(\Instance3.un1_r_Count_10lt11_0 ));
    InMux I__1421 (
            .O(N__6468),
            .I(N__6465));
    LocalMux I__1420 (
            .O(N__6465),
            .I(\Instance3.un1_r_Count_10lto11_1 ));
    InMux I__1419 (
            .O(N__6462),
            .I(N__6459));
    LocalMux I__1418 (
            .O(N__6459),
            .I(\Instance3.r_Count13_4 ));
    CascadeMux I__1417 (
            .O(N__6456),
            .I(N__6450));
    InMux I__1416 (
            .O(N__6455),
            .I(N__6445));
    InMux I__1415 (
            .O(N__6454),
            .I(N__6445));
    InMux I__1414 (
            .O(N__6453),
            .I(N__6442));
    InMux I__1413 (
            .O(N__6450),
            .I(N__6439));
    LocalMux I__1412 (
            .O(N__6445),
            .I(\Instance4.r_CountZ0Z_0 ));
    LocalMux I__1411 (
            .O(N__6442),
            .I(\Instance4.r_CountZ0Z_0 ));
    LocalMux I__1410 (
            .O(N__6439),
            .I(\Instance4.r_CountZ0Z_0 ));
    CascadeMux I__1409 (
            .O(N__6432),
            .I(\Instance4.r_Count13_8_0_cascade_ ));
    CascadeMux I__1408 (
            .O(N__6429),
            .I(N__6424));
    InMux I__1407 (
            .O(N__6428),
            .I(N__6421));
    InMux I__1406 (
            .O(N__6427),
            .I(N__6418));
    InMux I__1405 (
            .O(N__6424),
            .I(N__6415));
    LocalMux I__1404 (
            .O(N__6421),
            .I(\Instance4.r_CountZ0Z_5 ));
    LocalMux I__1403 (
            .O(N__6418),
            .I(\Instance4.r_CountZ0Z_5 ));
    LocalMux I__1402 (
            .O(N__6415),
            .I(\Instance4.r_CountZ0Z_5 ));
    InMux I__1401 (
            .O(N__6408),
            .I(N__6405));
    LocalMux I__1400 (
            .O(N__6405),
            .I(\Instance4.r_Count13_7 ));
    CascadeMux I__1399 (
            .O(N__6402),
            .I(\Instance4.r_Count13_13_cascade_ ));
    InMux I__1398 (
            .O(N__6399),
            .I(N__6396));
    LocalMux I__1397 (
            .O(N__6396),
            .I(N__6393));
    Odrv4 I__1396 (
            .O(N__6393),
            .I(\Instance4.r_Count13_12 ));
    CascadeMux I__1395 (
            .O(N__6390),
            .I(N__6385));
    InMux I__1394 (
            .O(N__6389),
            .I(N__6382));
    InMux I__1393 (
            .O(N__6388),
            .I(N__6377));
    InMux I__1392 (
            .O(N__6385),
            .I(N__6377));
    LocalMux I__1391 (
            .O(N__6382),
            .I(\Instance4.r_CountZ0Z_14 ));
    LocalMux I__1390 (
            .O(N__6377),
            .I(\Instance4.r_CountZ0Z_14 ));
    InMux I__1389 (
            .O(N__6372),
            .I(N__6367));
    InMux I__1388 (
            .O(N__6371),
            .I(N__6362));
    InMux I__1387 (
            .O(N__6370),
            .I(N__6362));
    LocalMux I__1386 (
            .O(N__6367),
            .I(\Instance4.r_CountZ0Z_17 ));
    LocalMux I__1385 (
            .O(N__6362),
            .I(\Instance4.r_CountZ0Z_17 ));
    InMux I__1384 (
            .O(N__6357),
            .I(N__6354));
    LocalMux I__1383 (
            .O(N__6354),
            .I(\Instance4.r_Count13_4 ));
    InMux I__1382 (
            .O(N__6351),
            .I(N__6346));
    InMux I__1381 (
            .O(N__6350),
            .I(N__6341));
    InMux I__1380 (
            .O(N__6349),
            .I(N__6341));
    LocalMux I__1379 (
            .O(N__6346),
            .I(\Instance4.r_CountZ0Z_11 ));
    LocalMux I__1378 (
            .O(N__6341),
            .I(\Instance4.r_CountZ0Z_11 ));
    CascadeMux I__1377 (
            .O(N__6336),
            .I(N__6331));
    InMux I__1376 (
            .O(N__6335),
            .I(N__6328));
    InMux I__1375 (
            .O(N__6334),
            .I(N__6323));
    InMux I__1374 (
            .O(N__6331),
            .I(N__6323));
    LocalMux I__1373 (
            .O(N__6328),
            .I(\Instance4.r_CountZ0Z_10 ));
    LocalMux I__1372 (
            .O(N__6323),
            .I(\Instance4.r_CountZ0Z_10 ));
    InMux I__1371 (
            .O(N__6318),
            .I(N__6313));
    InMux I__1370 (
            .O(N__6317),
            .I(N__6310));
    InMux I__1369 (
            .O(N__6316),
            .I(N__6307));
    LocalMux I__1368 (
            .O(N__6313),
            .I(\Instance4.r_CountZ0Z_9 ));
    LocalMux I__1367 (
            .O(N__6310),
            .I(\Instance4.r_CountZ0Z_9 ));
    LocalMux I__1366 (
            .O(N__6307),
            .I(\Instance4.r_CountZ0Z_9 ));
    InMux I__1365 (
            .O(N__6300),
            .I(N__6295));
    InMux I__1364 (
            .O(N__6299),
            .I(N__6292));
    InMux I__1363 (
            .O(N__6298),
            .I(N__6289));
    LocalMux I__1362 (
            .O(N__6295),
            .I(\Instance4.r_CountZ0Z_13 ));
    LocalMux I__1361 (
            .O(N__6292),
            .I(\Instance4.r_CountZ0Z_13 ));
    LocalMux I__1360 (
            .O(N__6289),
            .I(\Instance4.r_CountZ0Z_13 ));
    InMux I__1359 (
            .O(N__6282),
            .I(N__6277));
    InMux I__1358 (
            .O(N__6281),
            .I(N__6274));
    InMux I__1357 (
            .O(N__6280),
            .I(N__6271));
    LocalMux I__1356 (
            .O(N__6277),
            .I(\Instance4.r_CountZ0Z_12 ));
    LocalMux I__1355 (
            .O(N__6274),
            .I(\Instance4.r_CountZ0Z_12 ));
    LocalMux I__1354 (
            .O(N__6271),
            .I(\Instance4.r_CountZ0Z_12 ));
    CascadeMux I__1353 (
            .O(N__6264),
            .I(\Instance4.un1_r_Count_10lto11_1_cascade_ ));
    InMux I__1352 (
            .O(N__6261),
            .I(N__6258));
    LocalMux I__1351 (
            .O(N__6258),
            .I(\Instance4.un1_r_Count_10lt11_0 ));
    InMux I__1350 (
            .O(N__6255),
            .I(N__6249));
    InMux I__1349 (
            .O(N__6254),
            .I(N__6249));
    LocalMux I__1348 (
            .O(N__6249),
            .I(N__6246));
    Span4Mux_v I__1347 (
            .O(N__6246),
            .I(N__6243));
    Span4Mux_h I__1346 (
            .O(N__6243),
            .I(N__6240));
    Odrv4 I__1345 (
            .O(N__6240),
            .I(i_Switch_4_c));
    InMux I__1344 (
            .O(N__6237),
            .I(N__6231));
    InMux I__1343 (
            .O(N__6236),
            .I(N__6231));
    LocalMux I__1342 (
            .O(N__6231),
            .I(N__6228));
    Span4Mux_v I__1341 (
            .O(N__6228),
            .I(N__6223));
    InMux I__1340 (
            .O(N__6227),
            .I(N__6218));
    InMux I__1339 (
            .O(N__6226),
            .I(N__6218));
    Odrv4 I__1338 (
            .O(N__6223),
            .I(w_Switch_4));
    LocalMux I__1337 (
            .O(N__6218),
            .I(w_Switch_4));
    CascadeMux I__1336 (
            .O(N__6213),
            .I(\Instance4.un1_r_Count_10lt17_cascade_ ));
    InMux I__1335 (
            .O(N__6210),
            .I(N__6207));
    LocalMux I__1334 (
            .O(N__6207),
            .I(\Instance4.un1_r_Count_10lto17_1 ));
    IoInMux I__1333 (
            .O(N__6204),
            .I(N__6201));
    LocalMux I__1332 (
            .O(N__6201),
            .I(N__6198));
    Span12Mux_s1_v I__1331 (
            .O(N__6198),
            .I(N__6195));
    Odrv12 I__1330 (
            .O(N__6195),
            .I(\Instance4.r_Count12_i ));
    InMux I__1329 (
            .O(N__6192),
            .I(bfn_6_12_0_));
    InMux I__1328 (
            .O(N__6189),
            .I(N__6184));
    InMux I__1327 (
            .O(N__6188),
            .I(N__6181));
    InMux I__1326 (
            .O(N__6187),
            .I(N__6178));
    LocalMux I__1325 (
            .O(N__6184),
            .I(\Instance2.r_CountZ0Z_17 ));
    LocalMux I__1324 (
            .O(N__6181),
            .I(\Instance2.r_CountZ0Z_17 ));
    LocalMux I__1323 (
            .O(N__6178),
            .I(\Instance2.r_CountZ0Z_17 ));
    CascadeMux I__1322 (
            .O(N__6171),
            .I(N__6167));
    InMux I__1321 (
            .O(N__6170),
            .I(N__6162));
    InMux I__1320 (
            .O(N__6167),
            .I(N__6159));
    InMux I__1319 (
            .O(N__6166),
            .I(N__6154));
    InMux I__1318 (
            .O(N__6165),
            .I(N__6154));
    LocalMux I__1317 (
            .O(N__6162),
            .I(N__6149));
    LocalMux I__1316 (
            .O(N__6159),
            .I(N__6149));
    LocalMux I__1315 (
            .O(N__6154),
            .I(\Instance2.r_Count_0_0 ));
    Odrv4 I__1314 (
            .O(N__6149),
            .I(\Instance2.r_Count_0_0 ));
    InMux I__1313 (
            .O(N__6144),
            .I(N__6139));
    CascadeMux I__1312 (
            .O(N__6143),
            .I(N__6136));
    InMux I__1311 (
            .O(N__6142),
            .I(N__6133));
    LocalMux I__1310 (
            .O(N__6139),
            .I(N__6130));
    InMux I__1309 (
            .O(N__6136),
            .I(N__6127));
    LocalMux I__1308 (
            .O(N__6133),
            .I(\Instance2.r_Count_0_1 ));
    Odrv4 I__1307 (
            .O(N__6130),
            .I(\Instance2.r_Count_0_1 ));
    LocalMux I__1306 (
            .O(N__6127),
            .I(\Instance2.r_Count_0_1 ));
    SRMux I__1305 (
            .O(N__6120),
            .I(N__6111));
    SRMux I__1304 (
            .O(N__6119),
            .I(N__6111));
    SRMux I__1303 (
            .O(N__6118),
            .I(N__6111));
    GlobalMux I__1302 (
            .O(N__6111),
            .I(N__6108));
    gio2CtrlBuf I__1301 (
            .O(N__6108),
            .I(\Instance2.r_Count12_i_g ));
    InMux I__1300 (
            .O(N__6105),
            .I(N__6102));
    LocalMux I__1299 (
            .O(N__6102),
            .I(N__6099));
    Span4Mux_v I__1298 (
            .O(N__6099),
            .I(N__6095));
    InMux I__1297 (
            .O(N__6098),
            .I(N__6092));
    Odrv4 I__1296 (
            .O(N__6095),
            .I(CONSTANT_ONE_NET));
    LocalMux I__1295 (
            .O(N__6092),
            .I(CONSTANT_ONE_NET));
    IoInMux I__1294 (
            .O(N__6087),
            .I(N__6084));
    LocalMux I__1293 (
            .O(N__6084),
            .I(N__6081));
    Odrv12 I__1292 (
            .O(N__6081),
            .I(r_HexEncode_i_0_3));
    InMux I__1291 (
            .O(N__6078),
            .I(N__6073));
    InMux I__1290 (
            .O(N__6077),
            .I(N__6068));
    InMux I__1289 (
            .O(N__6076),
            .I(N__6068));
    LocalMux I__1288 (
            .O(N__6073),
            .I(N__6061));
    LocalMux I__1287 (
            .O(N__6068),
            .I(N__6061));
    InMux I__1286 (
            .O(N__6067),
            .I(N__6054));
    InMux I__1285 (
            .O(N__6066),
            .I(N__6054));
    Span4Mux_h I__1284 (
            .O(N__6061),
            .I(N__6051));
    InMux I__1283 (
            .O(N__6060),
            .I(N__6046));
    InMux I__1282 (
            .O(N__6059),
            .I(N__6046));
    LocalMux I__1281 (
            .O(N__6054),
            .I(N__6043));
    Span4Mux_h I__1280 (
            .O(N__6051),
            .I(N__6040));
    LocalMux I__1279 (
            .O(N__6046),
            .I(sevseglZ0Z_2));
    Odrv4 I__1278 (
            .O(N__6043),
            .I(sevseglZ0Z_2));
    Odrv4 I__1277 (
            .O(N__6040),
            .I(sevseglZ0Z_2));
    InMux I__1276 (
            .O(N__6033),
            .I(N__6025));
    InMux I__1275 (
            .O(N__6032),
            .I(N__6025));
    InMux I__1274 (
            .O(N__6031),
            .I(N__6022));
    CascadeMux I__1273 (
            .O(N__6030),
            .I(N__6019));
    LocalMux I__1272 (
            .O(N__6025),
            .I(N__6011));
    LocalMux I__1271 (
            .O(N__6022),
            .I(N__6011));
    InMux I__1270 (
            .O(N__6019),
            .I(N__6006));
    InMux I__1269 (
            .O(N__6018),
            .I(N__6006));
    InMux I__1268 (
            .O(N__6017),
            .I(N__6001));
    InMux I__1267 (
            .O(N__6016),
            .I(N__6001));
    Span4Mux_s3_v I__1266 (
            .O(N__6011),
            .I(N__5998));
    LocalMux I__1265 (
            .O(N__6006),
            .I(sevseglZ0Z_1));
    LocalMux I__1264 (
            .O(N__6001),
            .I(sevseglZ0Z_1));
    Odrv4 I__1263 (
            .O(N__5998),
            .I(sevseglZ0Z_1));
    CascadeMux I__1262 (
            .O(N__5991),
            .I(N__5986));
    CascadeMux I__1261 (
            .O(N__5990),
            .I(N__5983));
    CascadeMux I__1260 (
            .O(N__5989),
            .I(N__5980));
    InMux I__1259 (
            .O(N__5986),
            .I(N__5975));
    InMux I__1258 (
            .O(N__5983),
            .I(N__5975));
    InMux I__1257 (
            .O(N__5980),
            .I(N__5972));
    LocalMux I__1256 (
            .O(N__5975),
            .I(N__5964));
    LocalMux I__1255 (
            .O(N__5972),
            .I(N__5964));
    CascadeMux I__1254 (
            .O(N__5971),
            .I(N__5960));
    CascadeMux I__1253 (
            .O(N__5970),
            .I(N__5957));
    CascadeMux I__1252 (
            .O(N__5969),
            .I(N__5954));
    Span4Mux_h I__1251 (
            .O(N__5964),
            .I(N__5951));
    InMux I__1250 (
            .O(N__5963),
            .I(N__5946));
    InMux I__1249 (
            .O(N__5960),
            .I(N__5946));
    InMux I__1248 (
            .O(N__5957),
            .I(N__5941));
    InMux I__1247 (
            .O(N__5954),
            .I(N__5941));
    Odrv4 I__1246 (
            .O(N__5951),
            .I(sevseglZ0Z_3));
    LocalMux I__1245 (
            .O(N__5946),
            .I(sevseglZ0Z_3));
    LocalMux I__1244 (
            .O(N__5941),
            .I(sevseglZ0Z_3));
    InMux I__1243 (
            .O(N__5934),
            .I(N__5928));
    InMux I__1242 (
            .O(N__5933),
            .I(N__5928));
    LocalMux I__1241 (
            .O(N__5928),
            .I(N__5924));
    InMux I__1240 (
            .O(N__5927),
            .I(N__5921));
    Span4Mux_h I__1239 (
            .O(N__5924),
            .I(N__5916));
    LocalMux I__1238 (
            .O(N__5921),
            .I(N__5916));
    Span4Mux_h I__1237 (
            .O(N__5916),
            .I(N__5909));
    InMux I__1236 (
            .O(N__5915),
            .I(N__5904));
    InMux I__1235 (
            .O(N__5914),
            .I(N__5904));
    InMux I__1234 (
            .O(N__5913),
            .I(N__5899));
    InMux I__1233 (
            .O(N__5912),
            .I(N__5899));
    Odrv4 I__1232 (
            .O(N__5909),
            .I(sevseglZ0Z_0));
    LocalMux I__1231 (
            .O(N__5904),
            .I(sevseglZ0Z_0));
    LocalMux I__1230 (
            .O(N__5899),
            .I(sevseglZ0Z_0));
    IoInMux I__1229 (
            .O(N__5892),
            .I(N__5889));
    LocalMux I__1228 (
            .O(N__5889),
            .I(N__5886));
    Odrv4 I__1227 (
            .O(N__5886),
            .I(r_HexEncode_i_0_2));
    InMux I__1226 (
            .O(N__5883),
            .I(N__5878));
    InMux I__1225 (
            .O(N__5882),
            .I(N__5875));
    InMux I__1224 (
            .O(N__5881),
            .I(N__5872));
    LocalMux I__1223 (
            .O(N__5878),
            .I(\Instance4.r_CountZ0Z_1 ));
    LocalMux I__1222 (
            .O(N__5875),
            .I(\Instance4.r_CountZ0Z_1 ));
    LocalMux I__1221 (
            .O(N__5872),
            .I(\Instance4.r_CountZ0Z_1 ));
    InMux I__1220 (
            .O(N__5865),
            .I(N__5861));
    InMux I__1219 (
            .O(N__5864),
            .I(N__5858));
    LocalMux I__1218 (
            .O(N__5861),
            .I(\Instance4.r_CountZ0Z_2 ));
    LocalMux I__1217 (
            .O(N__5858),
            .I(\Instance4.r_CountZ0Z_2 ));
    CascadeMux I__1216 (
            .O(N__5853),
            .I(N__5849));
    InMux I__1215 (
            .O(N__5852),
            .I(N__5846));
    InMux I__1214 (
            .O(N__5849),
            .I(N__5843));
    LocalMux I__1213 (
            .O(N__5846),
            .I(\Instance4.r_CountZ0Z_3 ));
    LocalMux I__1212 (
            .O(N__5843),
            .I(\Instance4.r_CountZ0Z_3 ));
    InMux I__1211 (
            .O(N__5838),
            .I(N__5833));
    InMux I__1210 (
            .O(N__5837),
            .I(N__5828));
    InMux I__1209 (
            .O(N__5836),
            .I(N__5828));
    LocalMux I__1208 (
            .O(N__5833),
            .I(\Instance4.r_CountZ0Z_4 ));
    LocalMux I__1207 (
            .O(N__5828),
            .I(\Instance4.r_CountZ0Z_4 ));
    CascadeMux I__1206 (
            .O(N__5823),
            .I(N__5820));
    InMux I__1205 (
            .O(N__5820),
            .I(N__5815));
    InMux I__1204 (
            .O(N__5819),
            .I(N__5812));
    InMux I__1203 (
            .O(N__5818),
            .I(N__5809));
    LocalMux I__1202 (
            .O(N__5815),
            .I(\Instance4.r_CountZ0Z_7 ));
    LocalMux I__1201 (
            .O(N__5812),
            .I(\Instance4.r_CountZ0Z_7 ));
    LocalMux I__1200 (
            .O(N__5809),
            .I(\Instance4.r_CountZ0Z_7 ));
    InMux I__1199 (
            .O(N__5802),
            .I(N__5797));
    InMux I__1198 (
            .O(N__5801),
            .I(N__5792));
    InMux I__1197 (
            .O(N__5800),
            .I(N__5792));
    LocalMux I__1196 (
            .O(N__5797),
            .I(\Instance2.r_CountZ0Z_9 ));
    LocalMux I__1195 (
            .O(N__5792),
            .I(\Instance2.r_CountZ0Z_9 ));
    InMux I__1194 (
            .O(N__5787),
            .I(bfn_6_11_0_));
    InMux I__1193 (
            .O(N__5784),
            .I(N__5779));
    InMux I__1192 (
            .O(N__5783),
            .I(N__5776));
    InMux I__1191 (
            .O(N__5782),
            .I(N__5773));
    LocalMux I__1190 (
            .O(N__5779),
            .I(N__5770));
    LocalMux I__1189 (
            .O(N__5776),
            .I(\Instance2.r_CountZ0Z_10 ));
    LocalMux I__1188 (
            .O(N__5773),
            .I(\Instance2.r_CountZ0Z_10 ));
    Odrv4 I__1187 (
            .O(N__5770),
            .I(\Instance2.r_CountZ0Z_10 ));
    InMux I__1186 (
            .O(N__5763),
            .I(\Instance2.r_Count_2_cry_9 ));
    CascadeMux I__1185 (
            .O(N__5760),
            .I(N__5755));
    InMux I__1184 (
            .O(N__5759),
            .I(N__5752));
    InMux I__1183 (
            .O(N__5758),
            .I(N__5749));
    InMux I__1182 (
            .O(N__5755),
            .I(N__5746));
    LocalMux I__1181 (
            .O(N__5752),
            .I(\Instance2.r_CountZ0Z_11 ));
    LocalMux I__1180 (
            .O(N__5749),
            .I(\Instance2.r_CountZ0Z_11 ));
    LocalMux I__1179 (
            .O(N__5746),
            .I(\Instance2.r_CountZ0Z_11 ));
    InMux I__1178 (
            .O(N__5739),
            .I(\Instance2.r_Count_2_cry_10 ));
    InMux I__1177 (
            .O(N__5736),
            .I(N__5731));
    InMux I__1176 (
            .O(N__5735),
            .I(N__5728));
    InMux I__1175 (
            .O(N__5734),
            .I(N__5725));
    LocalMux I__1174 (
            .O(N__5731),
            .I(\Instance2.r_CountZ0Z_12 ));
    LocalMux I__1173 (
            .O(N__5728),
            .I(\Instance2.r_CountZ0Z_12 ));
    LocalMux I__1172 (
            .O(N__5725),
            .I(\Instance2.r_CountZ0Z_12 ));
    InMux I__1171 (
            .O(N__5718),
            .I(\Instance2.r_Count_2_cry_11 ));
    CascadeMux I__1170 (
            .O(N__5715),
            .I(N__5711));
    InMux I__1169 (
            .O(N__5714),
            .I(N__5707));
    InMux I__1168 (
            .O(N__5711),
            .I(N__5702));
    InMux I__1167 (
            .O(N__5710),
            .I(N__5702));
    LocalMux I__1166 (
            .O(N__5707),
            .I(\Instance2.r_CountZ0Z_13 ));
    LocalMux I__1165 (
            .O(N__5702),
            .I(\Instance2.r_CountZ0Z_13 ));
    InMux I__1164 (
            .O(N__5697),
            .I(\Instance2.r_Count_2_cry_12 ));
    CascadeMux I__1163 (
            .O(N__5694),
            .I(N__5689));
    InMux I__1162 (
            .O(N__5693),
            .I(N__5686));
    InMux I__1161 (
            .O(N__5692),
            .I(N__5683));
    InMux I__1160 (
            .O(N__5689),
            .I(N__5680));
    LocalMux I__1159 (
            .O(N__5686),
            .I(\Instance2.r_CountZ0Z_14 ));
    LocalMux I__1158 (
            .O(N__5683),
            .I(\Instance2.r_CountZ0Z_14 ));
    LocalMux I__1157 (
            .O(N__5680),
            .I(\Instance2.r_CountZ0Z_14 ));
    InMux I__1156 (
            .O(N__5673),
            .I(\Instance2.r_Count_2_cry_13 ));
    CascadeMux I__1155 (
            .O(N__5670),
            .I(N__5666));
    InMux I__1154 (
            .O(N__5669),
            .I(N__5662));
    InMux I__1153 (
            .O(N__5666),
            .I(N__5659));
    InMux I__1152 (
            .O(N__5665),
            .I(N__5656));
    LocalMux I__1151 (
            .O(N__5662),
            .I(\Instance2.r_CountZ0Z_15 ));
    LocalMux I__1150 (
            .O(N__5659),
            .I(\Instance2.r_CountZ0Z_15 ));
    LocalMux I__1149 (
            .O(N__5656),
            .I(\Instance2.r_CountZ0Z_15 ));
    InMux I__1148 (
            .O(N__5649),
            .I(\Instance2.r_Count_2_cry_14 ));
    InMux I__1147 (
            .O(N__5646),
            .I(N__5642));
    InMux I__1146 (
            .O(N__5645),
            .I(N__5638));
    LocalMux I__1145 (
            .O(N__5642),
            .I(N__5635));
    InMux I__1144 (
            .O(N__5641),
            .I(N__5632));
    LocalMux I__1143 (
            .O(N__5638),
            .I(\Instance2.r_CountZ0Z_16 ));
    Odrv4 I__1142 (
            .O(N__5635),
            .I(\Instance2.r_CountZ0Z_16 ));
    LocalMux I__1141 (
            .O(N__5632),
            .I(\Instance2.r_CountZ0Z_16 ));
    InMux I__1140 (
            .O(N__5625),
            .I(\Instance2.r_Count_2_cry_15 ));
    SRMux I__1139 (
            .O(N__5622),
            .I(N__5610));
    SRMux I__1138 (
            .O(N__5621),
            .I(N__5610));
    SRMux I__1137 (
            .O(N__5620),
            .I(N__5610));
    SRMux I__1136 (
            .O(N__5619),
            .I(N__5610));
    GlobalMux I__1135 (
            .O(N__5610),
            .I(N__5607));
    gio2CtrlBuf I__1134 (
            .O(N__5607),
            .I(\Instance4.r_Count12_i_g ));
    InMux I__1133 (
            .O(N__5604),
            .I(N__5600));
    InMux I__1132 (
            .O(N__5603),
            .I(N__5597));
    LocalMux I__1131 (
            .O(N__5600),
            .I(\Instance2.r_Count_0_2 ));
    LocalMux I__1130 (
            .O(N__5597),
            .I(\Instance2.r_Count_0_2 ));
    InMux I__1129 (
            .O(N__5592),
            .I(\Instance2.r_Count_2_cry_1 ));
    InMux I__1128 (
            .O(N__5589),
            .I(N__5586));
    LocalMux I__1127 (
            .O(N__5586),
            .I(N__5583));
    Span4Mux_h I__1126 (
            .O(N__5583),
            .I(N__5579));
    InMux I__1125 (
            .O(N__5582),
            .I(N__5576));
    Odrv4 I__1124 (
            .O(N__5579),
            .I(\Instance2.r_Count_0_3 ));
    LocalMux I__1123 (
            .O(N__5576),
            .I(\Instance2.r_Count_0_3 ));
    InMux I__1122 (
            .O(N__5571),
            .I(\Instance2.r_Count_2_cry_2 ));
    InMux I__1121 (
            .O(N__5568),
            .I(N__5563));
    InMux I__1120 (
            .O(N__5567),
            .I(N__5560));
    InMux I__1119 (
            .O(N__5566),
            .I(N__5557));
    LocalMux I__1118 (
            .O(N__5563),
            .I(N__5552));
    LocalMux I__1117 (
            .O(N__5560),
            .I(N__5552));
    LocalMux I__1116 (
            .O(N__5557),
            .I(\Instance2.r_CountZ0Z_4 ));
    Odrv4 I__1115 (
            .O(N__5552),
            .I(\Instance2.r_CountZ0Z_4 ));
    InMux I__1114 (
            .O(N__5547),
            .I(\Instance2.r_Count_2_cry_3 ));
    InMux I__1113 (
            .O(N__5544),
            .I(N__5539));
    InMux I__1112 (
            .O(N__5543),
            .I(N__5534));
    InMux I__1111 (
            .O(N__5542),
            .I(N__5534));
    LocalMux I__1110 (
            .O(N__5539),
            .I(\Instance2.r_CountZ0Z_5 ));
    LocalMux I__1109 (
            .O(N__5534),
            .I(\Instance2.r_CountZ0Z_5 ));
    InMux I__1108 (
            .O(N__5529),
            .I(\Instance2.r_Count_2_cry_4 ));
    InMux I__1107 (
            .O(N__5526),
            .I(N__5521));
    InMux I__1106 (
            .O(N__5525),
            .I(N__5518));
    InMux I__1105 (
            .O(N__5524),
            .I(N__5515));
    LocalMux I__1104 (
            .O(N__5521),
            .I(\Instance2.r_CountZ0Z_6 ));
    LocalMux I__1103 (
            .O(N__5518),
            .I(\Instance2.r_CountZ0Z_6 ));
    LocalMux I__1102 (
            .O(N__5515),
            .I(\Instance2.r_CountZ0Z_6 ));
    InMux I__1101 (
            .O(N__5508),
            .I(\Instance2.r_Count_2_cry_5 ));
    CascadeMux I__1100 (
            .O(N__5505),
            .I(N__5500));
    InMux I__1099 (
            .O(N__5504),
            .I(N__5497));
    InMux I__1098 (
            .O(N__5503),
            .I(N__5494));
    InMux I__1097 (
            .O(N__5500),
            .I(N__5491));
    LocalMux I__1096 (
            .O(N__5497),
            .I(\Instance2.r_CountZ0Z_7 ));
    LocalMux I__1095 (
            .O(N__5494),
            .I(\Instance2.r_CountZ0Z_7 ));
    LocalMux I__1094 (
            .O(N__5491),
            .I(\Instance2.r_CountZ0Z_7 ));
    InMux I__1093 (
            .O(N__5484),
            .I(\Instance2.r_Count_2_cry_6 ));
    InMux I__1092 (
            .O(N__5481),
            .I(N__5476));
    InMux I__1091 (
            .O(N__5480),
            .I(N__5471));
    InMux I__1090 (
            .O(N__5479),
            .I(N__5471));
    LocalMux I__1089 (
            .O(N__5476),
            .I(\Instance2.r_CountZ0Z_8 ));
    LocalMux I__1088 (
            .O(N__5471),
            .I(\Instance2.r_CountZ0Z_8 ));
    InMux I__1087 (
            .O(N__5466),
            .I(\Instance2.r_Count_2_cry_7 ));
    InMux I__1086 (
            .O(N__5463),
            .I(bfn_6_8_0_));
    InMux I__1085 (
            .O(N__5460),
            .I(\Instance4.r_Count_2_cry_9 ));
    InMux I__1084 (
            .O(N__5457),
            .I(\Instance4.r_Count_2_cry_10 ));
    InMux I__1083 (
            .O(N__5454),
            .I(\Instance4.r_Count_2_cry_11 ));
    InMux I__1082 (
            .O(N__5451),
            .I(\Instance4.r_Count_2_cry_12 ));
    InMux I__1081 (
            .O(N__5448),
            .I(\Instance4.r_Count_2_cry_13 ));
    InMux I__1080 (
            .O(N__5445),
            .I(\Instance4.r_Count_2_cry_14 ));
    InMux I__1079 (
            .O(N__5442),
            .I(\Instance4.r_Count_2_cry_15 ));
    InMux I__1078 (
            .O(N__5439),
            .I(bfn_6_9_0_));
    InMux I__1077 (
            .O(N__5436),
            .I(\Instance4.r_Count_2_cry_1 ));
    InMux I__1076 (
            .O(N__5433),
            .I(\Instance4.r_Count_2_cry_2 ));
    InMux I__1075 (
            .O(N__5430),
            .I(\Instance4.r_Count_2_cry_3 ));
    InMux I__1074 (
            .O(N__5427),
            .I(\Instance4.r_Count_2_cry_4 ));
    InMux I__1073 (
            .O(N__5424),
            .I(\Instance4.r_Count_2_cry_5 ));
    InMux I__1072 (
            .O(N__5421),
            .I(\Instance4.r_Count_2_cry_6 ));
    InMux I__1071 (
            .O(N__5418),
            .I(\Instance4.r_Count_2_cry_7 ));
    IoInMux I__1070 (
            .O(N__5415),
            .I(N__5412));
    LocalMux I__1069 (
            .O(N__5412),
            .I(N__5409));
    Odrv4 I__1068 (
            .O(N__5409),
            .I(r_HexEncode_i_0_4));
    CEMux I__1067 (
            .O(N__5406),
            .I(N__5401));
    CEMux I__1066 (
            .O(N__5405),
            .I(N__5397));
    CEMux I__1065 (
            .O(N__5404),
            .I(N__5394));
    LocalMux I__1064 (
            .O(N__5401),
            .I(N__5391));
    CEMux I__1063 (
            .O(N__5400),
            .I(N__5388));
    LocalMux I__1062 (
            .O(N__5397),
            .I(N__5383));
    LocalMux I__1061 (
            .O(N__5394),
            .I(N__5383));
    Span4Mux_v I__1060 (
            .O(N__5391),
            .I(N__5380));
    LocalMux I__1059 (
            .O(N__5388),
            .I(N__5377));
    Span4Mux_h I__1058 (
            .O(N__5383),
            .I(N__5374));
    Span4Mux_h I__1057 (
            .O(N__5380),
            .I(N__5369));
    Span4Mux_h I__1056 (
            .O(N__5377),
            .I(N__5369));
    Odrv4 I__1055 (
            .O(N__5374),
            .I(\alogicunit.N_35 ));
    Odrv4 I__1054 (
            .O(N__5369),
            .I(\alogicunit.N_35 ));
    InMux I__1053 (
            .O(N__5364),
            .I(N__5358));
    InMux I__1052 (
            .O(N__5363),
            .I(N__5358));
    LocalMux I__1051 (
            .O(N__5358),
            .I(N__5352));
    InMux I__1050 (
            .O(N__5357),
            .I(N__5347));
    InMux I__1049 (
            .O(N__5356),
            .I(N__5347));
    InMux I__1048 (
            .O(N__5355),
            .I(N__5344));
    Odrv4 I__1047 (
            .O(N__5352),
            .I(\alogicunit.result24_iZ0 ));
    LocalMux I__1046 (
            .O(N__5347),
            .I(\alogicunit.result24_iZ0 ));
    LocalMux I__1045 (
            .O(N__5344),
            .I(\alogicunit.result24_iZ0 ));
    InMux I__1044 (
            .O(N__5337),
            .I(N__5332));
    CascadeMux I__1043 (
            .O(N__5336),
            .I(N__5329));
    CascadeMux I__1042 (
            .O(N__5335),
            .I(N__5324));
    LocalMux I__1041 (
            .O(N__5332),
            .I(N__5316));
    InMux I__1040 (
            .O(N__5329),
            .I(N__5312));
    InMux I__1039 (
            .O(N__5328),
            .I(N__5307));
    InMux I__1038 (
            .O(N__5327),
            .I(N__5307));
    InMux I__1037 (
            .O(N__5324),
            .I(N__5304));
    CascadeMux I__1036 (
            .O(N__5323),
            .I(N__5298));
    InMux I__1035 (
            .O(N__5322),
            .I(N__5291));
    InMux I__1034 (
            .O(N__5321),
            .I(N__5284));
    InMux I__1033 (
            .O(N__5320),
            .I(N__5284));
    InMux I__1032 (
            .O(N__5319),
            .I(N__5284));
    Span4Mux_h I__1031 (
            .O(N__5316),
            .I(N__5281));
    InMux I__1030 (
            .O(N__5315),
            .I(N__5278));
    LocalMux I__1029 (
            .O(N__5312),
            .I(N__5271));
    LocalMux I__1028 (
            .O(N__5307),
            .I(N__5271));
    LocalMux I__1027 (
            .O(N__5304),
            .I(N__5271));
    InMux I__1026 (
            .O(N__5303),
            .I(N__5260));
    InMux I__1025 (
            .O(N__5302),
            .I(N__5260));
    InMux I__1024 (
            .O(N__5301),
            .I(N__5260));
    InMux I__1023 (
            .O(N__5298),
            .I(N__5260));
    InMux I__1022 (
            .O(N__5297),
            .I(N__5260));
    InMux I__1021 (
            .O(N__5296),
            .I(N__5257));
    InMux I__1020 (
            .O(N__5295),
            .I(N__5252));
    InMux I__1019 (
            .O(N__5294),
            .I(N__5252));
    LocalMux I__1018 (
            .O(N__5291),
            .I(current_state_0));
    LocalMux I__1017 (
            .O(N__5284),
            .I(current_state_0));
    Odrv4 I__1016 (
            .O(N__5281),
            .I(current_state_0));
    LocalMux I__1015 (
            .O(N__5278),
            .I(current_state_0));
    Odrv4 I__1014 (
            .O(N__5271),
            .I(current_state_0));
    LocalMux I__1013 (
            .O(N__5260),
            .I(current_state_0));
    LocalMux I__1012 (
            .O(N__5257),
            .I(current_state_0));
    LocalMux I__1011 (
            .O(N__5252),
            .I(current_state_0));
    CascadeMux I__1010 (
            .O(N__5235),
            .I(N__5231));
    CascadeMux I__1009 (
            .O(N__5234),
            .I(N__5228));
    InMux I__1008 (
            .O(N__5231),
            .I(N__5217));
    InMux I__1007 (
            .O(N__5228),
            .I(N__5217));
    InMux I__1006 (
            .O(N__5227),
            .I(N__5214));
    InMux I__1005 (
            .O(N__5226),
            .I(N__5211));
    CascadeMux I__1004 (
            .O(N__5225),
            .I(N__5203));
    CascadeMux I__1003 (
            .O(N__5224),
            .I(N__5197));
    InMux I__1002 (
            .O(N__5223),
            .I(N__5194));
    InMux I__1001 (
            .O(N__5222),
            .I(N__5191));
    LocalMux I__1000 (
            .O(N__5217),
            .I(N__5186));
    LocalMux I__999 (
            .O(N__5214),
            .I(N__5186));
    LocalMux I__998 (
            .O(N__5211),
            .I(N__5183));
    InMux I__997 (
            .O(N__5210),
            .I(N__5170));
    InMux I__996 (
            .O(N__5209),
            .I(N__5170));
    InMux I__995 (
            .O(N__5208),
            .I(N__5170));
    InMux I__994 (
            .O(N__5207),
            .I(N__5170));
    InMux I__993 (
            .O(N__5206),
            .I(N__5170));
    InMux I__992 (
            .O(N__5203),
            .I(N__5170));
    InMux I__991 (
            .O(N__5202),
            .I(N__5161));
    InMux I__990 (
            .O(N__5201),
            .I(N__5161));
    InMux I__989 (
            .O(N__5200),
            .I(N__5161));
    InMux I__988 (
            .O(N__5197),
            .I(N__5161));
    LocalMux I__987 (
            .O(N__5194),
            .I(current_state_1));
    LocalMux I__986 (
            .O(N__5191),
            .I(current_state_1));
    Odrv4 I__985 (
            .O(N__5186),
            .I(current_state_1));
    Odrv4 I__984 (
            .O(N__5183),
            .I(current_state_1));
    LocalMux I__983 (
            .O(N__5170),
            .I(current_state_1));
    LocalMux I__982 (
            .O(N__5161),
            .I(current_state_1));
    InMux I__981 (
            .O(N__5148),
            .I(N__5134));
    InMux I__980 (
            .O(N__5147),
            .I(N__5134));
    InMux I__979 (
            .O(N__5146),
            .I(N__5134));
    InMux I__978 (
            .O(N__5145),
            .I(N__5127));
    InMux I__977 (
            .O(N__5144),
            .I(N__5122));
    InMux I__976 (
            .O(N__5143),
            .I(N__5122));
    InMux I__975 (
            .O(N__5142),
            .I(N__5119));
    CascadeMux I__974 (
            .O(N__5141),
            .I(N__5115));
    LocalMux I__973 (
            .O(N__5134),
            .I(N__5112));
    CascadeMux I__972 (
            .O(N__5133),
            .I(N__5108));
    CascadeMux I__971 (
            .O(N__5132),
            .I(N__5103));
    InMux I__970 (
            .O(N__5131),
            .I(N__5097));
    InMux I__969 (
            .O(N__5130),
            .I(N__5094));
    LocalMux I__968 (
            .O(N__5127),
            .I(N__5089));
    LocalMux I__967 (
            .O(N__5122),
            .I(N__5089));
    LocalMux I__966 (
            .O(N__5119),
            .I(N__5086));
    InMux I__965 (
            .O(N__5118),
            .I(N__5081));
    InMux I__964 (
            .O(N__5115),
            .I(N__5081));
    Span4Mux_v I__963 (
            .O(N__5112),
            .I(N__5078));
    InMux I__962 (
            .O(N__5111),
            .I(N__5067));
    InMux I__961 (
            .O(N__5108),
            .I(N__5067));
    InMux I__960 (
            .O(N__5107),
            .I(N__5067));
    InMux I__959 (
            .O(N__5106),
            .I(N__5067));
    InMux I__958 (
            .O(N__5103),
            .I(N__5067));
    InMux I__957 (
            .O(N__5102),
            .I(N__5064));
    InMux I__956 (
            .O(N__5101),
            .I(N__5059));
    InMux I__955 (
            .O(N__5100),
            .I(N__5059));
    LocalMux I__954 (
            .O(N__5097),
            .I(current_state_2));
    LocalMux I__953 (
            .O(N__5094),
            .I(current_state_2));
    Odrv4 I__952 (
            .O(N__5089),
            .I(current_state_2));
    Odrv4 I__951 (
            .O(N__5086),
            .I(current_state_2));
    LocalMux I__950 (
            .O(N__5081),
            .I(current_state_2));
    Odrv4 I__949 (
            .O(N__5078),
            .I(current_state_2));
    LocalMux I__948 (
            .O(N__5067),
            .I(current_state_2));
    LocalMux I__947 (
            .O(N__5064),
            .I(current_state_2));
    LocalMux I__946 (
            .O(N__5059),
            .I(current_state_2));
    InMux I__945 (
            .O(N__5040),
            .I(N__5034));
    InMux I__944 (
            .O(N__5039),
            .I(N__5029));
    InMux I__943 (
            .O(N__5038),
            .I(N__5029));
    InMux I__942 (
            .O(N__5037),
            .I(N__5026));
    LocalMux I__941 (
            .O(N__5034),
            .I(N__5013));
    LocalMux I__940 (
            .O(N__5029),
            .I(N__5013));
    LocalMux I__939 (
            .O(N__5026),
            .I(N__5010));
    InMux I__938 (
            .O(N__5025),
            .I(N__5005));
    InMux I__937 (
            .O(N__5024),
            .I(N__5005));
    InMux I__936 (
            .O(N__5023),
            .I(N__4992));
    InMux I__935 (
            .O(N__5022),
            .I(N__4992));
    InMux I__934 (
            .O(N__5021),
            .I(N__4992));
    InMux I__933 (
            .O(N__5020),
            .I(N__4992));
    InMux I__932 (
            .O(N__5019),
            .I(N__4992));
    InMux I__931 (
            .O(N__5018),
            .I(N__4992));
    Span4Mux_v I__930 (
            .O(N__5013),
            .I(N__4979));
    Span4Mux_h I__929 (
            .O(N__5010),
            .I(N__4979));
    LocalMux I__928 (
            .O(N__5005),
            .I(N__4979));
    LocalMux I__927 (
            .O(N__4992),
            .I(N__4979));
    InMux I__926 (
            .O(N__4991),
            .I(N__4970));
    InMux I__925 (
            .O(N__4990),
            .I(N__4970));
    InMux I__924 (
            .O(N__4989),
            .I(N__4970));
    InMux I__923 (
            .O(N__4988),
            .I(N__4970));
    Odrv4 I__922 (
            .O(N__4979),
            .I(current_state_3));
    LocalMux I__921 (
            .O(N__4970),
            .I(current_state_3));
    CEMux I__920 (
            .O(N__4965),
            .I(N__4960));
    CascadeMux I__919 (
            .O(N__4964),
            .I(N__4956));
    InMux I__918 (
            .O(N__4963),
            .I(N__4952));
    LocalMux I__917 (
            .O(N__4960),
            .I(N__4949));
    InMux I__916 (
            .O(N__4959),
            .I(N__4946));
    InMux I__915 (
            .O(N__4956),
            .I(N__4941));
    InMux I__914 (
            .O(N__4955),
            .I(N__4941));
    LocalMux I__913 (
            .O(N__4952),
            .I(N__4938));
    Span4Mux_s2_v I__912 (
            .O(N__4949),
            .I(N__4931));
    LocalMux I__911 (
            .O(N__4946),
            .I(N__4931));
    LocalMux I__910 (
            .O(N__4941),
            .I(N__4931));
    Odrv4 I__909 (
            .O(N__4938),
            .I(clickZ0Z1));
    Odrv4 I__908 (
            .O(N__4931),
            .I(clickZ0Z1));
    InMux I__907 (
            .O(N__4926),
            .I(N__4923));
    LocalMux I__906 (
            .O(N__4923),
            .I(N__4920));
    Odrv12 I__905 (
            .O(N__4920),
            .I(\Instance2.un1_r_Count_10lto17_1 ));
    InMux I__904 (
            .O(N__4917),
            .I(N__4912));
    InMux I__903 (
            .O(N__4916),
            .I(N__4909));
    InMux I__902 (
            .O(N__4915),
            .I(N__4906));
    LocalMux I__901 (
            .O(N__4912),
            .I(N__4903));
    LocalMux I__900 (
            .O(N__4909),
            .I(N__4898));
    LocalMux I__899 (
            .O(N__4906),
            .I(N__4895));
    Span12Mux_s4_h I__898 (
            .O(N__4903),
            .I(N__4892));
    InMux I__897 (
            .O(N__4902),
            .I(N__4887));
    InMux I__896 (
            .O(N__4901),
            .I(N__4887));
    Odrv4 I__895 (
            .O(N__4898),
            .I(w_Switch_2));
    Odrv12 I__894 (
            .O(N__4895),
            .I(w_Switch_2));
    Odrv12 I__893 (
            .O(N__4892),
            .I(w_Switch_2));
    LocalMux I__892 (
            .O(N__4887),
            .I(w_Switch_2));
    CascadeMux I__891 (
            .O(N__4878),
            .I(N__4875));
    InMux I__890 (
            .O(N__4875),
            .I(N__4872));
    LocalMux I__889 (
            .O(N__4872),
            .I(N__4868));
    InMux I__888 (
            .O(N__4871),
            .I(N__4865));
    Span4Mux_s3_v I__887 (
            .O(N__4868),
            .I(N__4862));
    LocalMux I__886 (
            .O(N__4865),
            .I(N__4859));
    Sp12to4 I__885 (
            .O(N__4862),
            .I(N__4854));
    Sp12to4 I__884 (
            .O(N__4859),
            .I(N__4854));
    Span12Mux_v I__883 (
            .O(N__4854),
            .I(N__4851));
    Odrv12 I__882 (
            .O(N__4851),
            .I(i_Switch_2_c));
    InMux I__881 (
            .O(N__4848),
            .I(N__4845));
    LocalMux I__880 (
            .O(N__4845),
            .I(N__4842));
    Odrv12 I__879 (
            .O(N__4842),
            .I(\Instance2.un1_r_Count_10lt17 ));
    IoInMux I__878 (
            .O(N__4839),
            .I(N__4836));
    LocalMux I__877 (
            .O(N__4836),
            .I(\Instance2.r_Count12_i ));
    InMux I__876 (
            .O(N__4833),
            .I(N__4830));
    LocalMux I__875 (
            .O(N__4830),
            .I(N__4826));
    InMux I__874 (
            .O(N__4829),
            .I(N__4823));
    Odrv12 I__873 (
            .O(N__4826),
            .I(r_SwitchZ0Z_2));
    LocalMux I__872 (
            .O(N__4823),
            .I(r_SwitchZ0Z_2));
    InMux I__871 (
            .O(N__4818),
            .I(N__4815));
    LocalMux I__870 (
            .O(N__4815),
            .I(r_SwitchZ0Z_4));
    CascadeMux I__869 (
            .O(N__4812),
            .I(\Instance2.click14_sn_cascade_ ));
    InMux I__868 (
            .O(N__4809),
            .I(N__4802));
    InMux I__867 (
            .O(N__4808),
            .I(N__4797));
    InMux I__866 (
            .O(N__4807),
            .I(N__4797));
    InMux I__865 (
            .O(N__4806),
            .I(N__4794));
    CascadeMux I__864 (
            .O(N__4805),
            .I(N__4791));
    LocalMux I__863 (
            .O(N__4802),
            .I(N__4782));
    LocalMux I__862 (
            .O(N__4797),
            .I(N__4782));
    LocalMux I__861 (
            .O(N__4794),
            .I(N__4782));
    InMux I__860 (
            .O(N__4791),
            .I(N__4774));
    InMux I__859 (
            .O(N__4790),
            .I(N__4774));
    InMux I__858 (
            .O(N__4789),
            .I(N__4774));
    Span4Mux_v I__857 (
            .O(N__4782),
            .I(N__4771));
    InMux I__856 (
            .O(N__4781),
            .I(N__4768));
    LocalMux I__855 (
            .O(N__4774),
            .I(un1_click13_1_sn));
    Odrv4 I__854 (
            .O(N__4771),
            .I(un1_click13_1_sn));
    LocalMux I__853 (
            .O(N__4768),
            .I(un1_click13_1_sn));
    InMux I__852 (
            .O(N__4761),
            .I(N__4757));
    InMux I__851 (
            .O(N__4760),
            .I(N__4754));
    LocalMux I__850 (
            .O(N__4757),
            .I(N__4751));
    LocalMux I__849 (
            .O(N__4754),
            .I(Instance2_un1_click13_3_1));
    Odrv12 I__848 (
            .O(N__4751),
            .I(Instance2_un1_click13_3_1));
    InMux I__847 (
            .O(N__4746),
            .I(N__4743));
    LocalMux I__846 (
            .O(N__4743),
            .I(\alogicunit.result_RNO_0Z0Z_4 ));
    CascadeMux I__845 (
            .O(N__4740),
            .I(N__4737));
    InMux I__844 (
            .O(N__4737),
            .I(N__4734));
    LocalMux I__843 (
            .O(N__4734),
            .I(N__4731));
    Span4Mux_s2_h I__842 (
            .O(N__4731),
            .I(N__4728));
    Odrv4 I__841 (
            .O(N__4728),
            .I(left_0));
    InMux I__840 (
            .O(N__4725),
            .I(N__4719));
    InMux I__839 (
            .O(N__4724),
            .I(N__4719));
    LocalMux I__838 (
            .O(N__4719),
            .I(\alogicunit.N_50 ));
    InMux I__837 (
            .O(N__4716),
            .I(N__4713));
    LocalMux I__836 (
            .O(N__4713),
            .I(\alogicunit.result_RNO_0Z0Z_6 ));
    InMux I__835 (
            .O(N__4710),
            .I(N__4707));
    LocalMux I__834 (
            .O(N__4707),
            .I(N__4704));
    Span4Mux_s2_h I__833 (
            .O(N__4704),
            .I(N__4701));
    Odrv4 I__832 (
            .O(N__4701),
            .I(left_2));
    InMux I__831 (
            .O(N__4698),
            .I(N__4694));
    InMux I__830 (
            .O(N__4697),
            .I(N__4691));
    LocalMux I__829 (
            .O(N__4694),
            .I(\alogicunit.un1_a_1_cry_1_c_invZ0 ));
    LocalMux I__828 (
            .O(N__4691),
            .I(\alogicunit.un1_a_1_cry_1_c_invZ0 ));
    InMux I__827 (
            .O(N__4686),
            .I(N__4680));
    InMux I__826 (
            .O(N__4685),
            .I(N__4680));
    LocalMux I__825 (
            .O(N__4680),
            .I(\alogicunit.N_102 ));
    InMux I__824 (
            .O(N__4677),
            .I(N__4674));
    LocalMux I__823 (
            .O(N__4674),
            .I(\Instance2.r_Count13_12 ));
    CascadeMux I__822 (
            .O(N__4671),
            .I(\Instance2.r_Count13_13_cascade_ ));
    InMux I__821 (
            .O(N__4668),
            .I(N__4665));
    LocalMux I__820 (
            .O(N__4665),
            .I(\Instance2.un1_r_Count_10lto11_1 ));
    CascadeMux I__819 (
            .O(N__4662),
            .I(N__4659));
    InMux I__818 (
            .O(N__4659),
            .I(N__4656));
    LocalMux I__817 (
            .O(N__4656),
            .I(\Instance2.r_Count13_10 ));
    InMux I__816 (
            .O(N__4653),
            .I(N__4650));
    LocalMux I__815 (
            .O(N__4650),
            .I(\Instance2.r_Count13_7 ));
    CascadeMux I__814 (
            .O(N__4647),
            .I(N__4644));
    InMux I__813 (
            .O(N__4644),
            .I(N__4638));
    InMux I__812 (
            .O(N__4643),
            .I(N__4638));
    LocalMux I__811 (
            .O(N__4638),
            .I(\alogicunit.N_90 ));
    InMux I__810 (
            .O(N__4635),
            .I(N__4632));
    LocalMux I__809 (
            .O(N__4632),
            .I(\Instance2.r_Count13_4 ));
    CEMux I__808 (
            .O(N__4629),
            .I(N__4626));
    LocalMux I__807 (
            .O(N__4626),
            .I(N__4617));
    InMux I__806 (
            .O(N__4625),
            .I(N__4614));
    InMux I__805 (
            .O(N__4624),
            .I(N__4607));
    InMux I__804 (
            .O(N__4623),
            .I(N__4607));
    InMux I__803 (
            .O(N__4622),
            .I(N__4607));
    InMux I__802 (
            .O(N__4621),
            .I(N__4599));
    InMux I__801 (
            .O(N__4620),
            .I(N__4599));
    Span4Mux_h I__800 (
            .O(N__4617),
            .I(N__4594));
    LocalMux I__799 (
            .O(N__4614),
            .I(N__4594));
    LocalMux I__798 (
            .O(N__4607),
            .I(N__4591));
    InMux I__797 (
            .O(N__4606),
            .I(N__4588));
    InMux I__796 (
            .O(N__4605),
            .I(N__4583));
    InMux I__795 (
            .O(N__4604),
            .I(N__4583));
    LocalMux I__794 (
            .O(N__4599),
            .I(N__4575));
    Span4Mux_v I__793 (
            .O(N__4594),
            .I(N__4570));
    Span4Mux_v I__792 (
            .O(N__4591),
            .I(N__4570));
    LocalMux I__791 (
            .O(N__4588),
            .I(N__4567));
    LocalMux I__790 (
            .O(N__4583),
            .I(N__4564));
    InMux I__789 (
            .O(N__4582),
            .I(N__4557));
    InMux I__788 (
            .O(N__4581),
            .I(N__4557));
    InMux I__787 (
            .O(N__4580),
            .I(N__4557));
    InMux I__786 (
            .O(N__4579),
            .I(N__4552));
    InMux I__785 (
            .O(N__4578),
            .I(N__4552));
    Odrv4 I__784 (
            .O(N__4575),
            .I(click13));
    Odrv4 I__783 (
            .O(N__4570),
            .I(click13));
    Odrv12 I__782 (
            .O(N__4567),
            .I(click13));
    Odrv4 I__781 (
            .O(N__4564),
            .I(click13));
    LocalMux I__780 (
            .O(N__4557),
            .I(click13));
    LocalMux I__779 (
            .O(N__4552),
            .I(click13));
    InMux I__778 (
            .O(N__4539),
            .I(N__4535));
    InMux I__777 (
            .O(N__4538),
            .I(N__4532));
    LocalMux I__776 (
            .O(N__4535),
            .I(\alogicunit.N_49 ));
    LocalMux I__775 (
            .O(N__4532),
            .I(\alogicunit.N_49 ));
    InMux I__774 (
            .O(N__4527),
            .I(N__4524));
    LocalMux I__773 (
            .O(N__4524),
            .I(N__4521));
    Span4Mux_s3_h I__772 (
            .O(N__4521),
            .I(N__4517));
    InMux I__771 (
            .O(N__4520),
            .I(N__4514));
    Odrv4 I__770 (
            .O(N__4517),
            .I(N_28));
    LocalMux I__769 (
            .O(N__4514),
            .I(N_28));
    InMux I__768 (
            .O(N__4509),
            .I(N__4503));
    InMux I__767 (
            .O(N__4508),
            .I(N__4503));
    LocalMux I__766 (
            .O(N__4503),
            .I(N__4500));
    Span4Mux_s3_h I__765 (
            .O(N__4500),
            .I(N__4497));
    Odrv4 I__764 (
            .O(N__4497),
            .I(\alogicunit.N_41 ));
    CascadeMux I__763 (
            .O(N__4494),
            .I(\alogicunit.N_41_cascade_ ));
    CascadeMux I__762 (
            .O(N__4491),
            .I(N__4487));
    CascadeMux I__761 (
            .O(N__4490),
            .I(N__4484));
    InMux I__760 (
            .O(N__4487),
            .I(N__4481));
    InMux I__759 (
            .O(N__4484),
            .I(N__4478));
    LocalMux I__758 (
            .O(N__4481),
            .I(N__4475));
    LocalMux I__757 (
            .O(N__4478),
            .I(N__4472));
    Span4Mux_s3_h I__756 (
            .O(N__4475),
            .I(N__4469));
    Span4Mux_v I__755 (
            .O(N__4472),
            .I(N__4466));
    Odrv4 I__754 (
            .O(N__4469),
            .I(track_RNI9MAL_0_1));
    Odrv4 I__753 (
            .O(N__4466),
            .I(track_RNI9MAL_0_1));
    CascadeMux I__752 (
            .O(N__4461),
            .I(N__4456));
    InMux I__751 (
            .O(N__4460),
            .I(N__4450));
    InMux I__750 (
            .O(N__4459),
            .I(N__4447));
    InMux I__749 (
            .O(N__4456),
            .I(N__4442));
    InMux I__748 (
            .O(N__4455),
            .I(N__4442));
    InMux I__747 (
            .O(N__4454),
            .I(N__4439));
    InMux I__746 (
            .O(N__4453),
            .I(N__4435));
    LocalMux I__745 (
            .O(N__4450),
            .I(N__4432));
    LocalMux I__744 (
            .O(N__4447),
            .I(N__4429));
    LocalMux I__743 (
            .O(N__4442),
            .I(N__4426));
    LocalMux I__742 (
            .O(N__4439),
            .I(N__4423));
    CascadeMux I__741 (
            .O(N__4438),
            .I(N__4420));
    LocalMux I__740 (
            .O(N__4435),
            .I(N__4415));
    Span4Mux_v I__739 (
            .O(N__4432),
            .I(N__4410));
    Span4Mux_v I__738 (
            .O(N__4429),
            .I(N__4410));
    Span4Mux_h I__737 (
            .O(N__4426),
            .I(N__4405));
    Span4Mux_s3_h I__736 (
            .O(N__4423),
            .I(N__4405));
    InMux I__735 (
            .O(N__4420),
            .I(N__4398));
    InMux I__734 (
            .O(N__4419),
            .I(N__4398));
    InMux I__733 (
            .O(N__4418),
            .I(N__4398));
    Odrv12 I__732 (
            .O(N__4415),
            .I(r_CountZ0Z_1));
    Odrv4 I__731 (
            .O(N__4410),
            .I(r_CountZ0Z_1));
    Odrv4 I__730 (
            .O(N__4405),
            .I(r_CountZ0Z_1));
    LocalMux I__729 (
            .O(N__4398),
            .I(r_CountZ0Z_1));
    InMux I__728 (
            .O(N__4389),
            .I(N__4377));
    InMux I__727 (
            .O(N__4388),
            .I(N__4377));
    InMux I__726 (
            .O(N__4387),
            .I(N__4377));
    InMux I__725 (
            .O(N__4386),
            .I(N__4372));
    InMux I__724 (
            .O(N__4385),
            .I(N__4372));
    InMux I__723 (
            .O(N__4384),
            .I(N__4369));
    LocalMux I__722 (
            .O(N__4377),
            .I(N__4366));
    LocalMux I__721 (
            .O(N__4372),
            .I(N__4363));
    LocalMux I__720 (
            .O(N__4369),
            .I(N__4356));
    Span4Mux_s3_h I__719 (
            .O(N__4366),
            .I(N__4353));
    Span4Mux_s3_h I__718 (
            .O(N__4363),
            .I(N__4350));
    InMux I__717 (
            .O(N__4362),
            .I(N__4341));
    InMux I__716 (
            .O(N__4361),
            .I(N__4341));
    InMux I__715 (
            .O(N__4360),
            .I(N__4341));
    InMux I__714 (
            .O(N__4359),
            .I(N__4341));
    Odrv12 I__713 (
            .O(N__4356),
            .I(r_CountZ0Z_0));
    Odrv4 I__712 (
            .O(N__4353),
            .I(r_CountZ0Z_0));
    Odrv4 I__711 (
            .O(N__4350),
            .I(r_CountZ0Z_0));
    LocalMux I__710 (
            .O(N__4341),
            .I(r_CountZ0Z_0));
    InMux I__709 (
            .O(N__4332),
            .I(N__4328));
    InMux I__708 (
            .O(N__4331),
            .I(N__4324));
    LocalMux I__707 (
            .O(N__4328),
            .I(N__4318));
    InMux I__706 (
            .O(N__4327),
            .I(N__4315));
    LocalMux I__705 (
            .O(N__4324),
            .I(N__4312));
    InMux I__704 (
            .O(N__4323),
            .I(N__4307));
    InMux I__703 (
            .O(N__4322),
            .I(N__4307));
    InMux I__702 (
            .O(N__4321),
            .I(N__4304));
    Span4Mux_h I__701 (
            .O(N__4318),
            .I(N__4301));
    LocalMux I__700 (
            .O(N__4315),
            .I(N__4298));
    Span4Mux_s3_h I__699 (
            .O(N__4312),
            .I(N__4295));
    LocalMux I__698 (
            .O(N__4307),
            .I(N__4292));
    LocalMux I__697 (
            .O(N__4304),
            .I(r_CountZ0Z_2));
    Odrv4 I__696 (
            .O(N__4301),
            .I(r_CountZ0Z_2));
    Odrv4 I__695 (
            .O(N__4298),
            .I(r_CountZ0Z_2));
    Odrv4 I__694 (
            .O(N__4295),
            .I(r_CountZ0Z_2));
    Odrv12 I__693 (
            .O(N__4292),
            .I(r_CountZ0Z_2));
    CascadeMux I__692 (
            .O(N__4281),
            .I(\Instance2.r_Count13_8_0_cascade_ ));
    CascadeMux I__691 (
            .O(N__4278),
            .I(\Instance2.un1_r_Count_10lt11_0_cascade_ ));
    InMux I__690 (
            .O(N__4275),
            .I(N__4272));
    LocalMux I__689 (
            .O(N__4272),
            .I(N__4269));
    Odrv4 I__688 (
            .O(N__4269),
            .I(sevsegr_RNO_0Z0Z_1));
    InMux I__687 (
            .O(N__4266),
            .I(N__4263));
    LocalMux I__686 (
            .O(N__4263),
            .I(r_SwitchZ0Z_3));
    CascadeMux I__685 (
            .O(N__4260),
            .I(N__4257));
    InMux I__684 (
            .O(N__4257),
            .I(N__4254));
    LocalMux I__683 (
            .O(N__4254),
            .I(\alogicunit.m26_l_fxZ0 ));
    InMux I__682 (
            .O(N__4251),
            .I(N__4248));
    LocalMux I__681 (
            .O(N__4248),
            .I(N__4245));
    Odrv4 I__680 (
            .O(N__4245),
            .I(sevsegl_RNO_0Z0Z_1));
    CascadeMux I__679 (
            .O(N__4242),
            .I(N__4239));
    InMux I__678 (
            .O(N__4239),
            .I(N__4235));
    CascadeMux I__677 (
            .O(N__4238),
            .I(N__4232));
    LocalMux I__676 (
            .O(N__4235),
            .I(N__4227));
    InMux I__675 (
            .O(N__4232),
            .I(N__4224));
    CascadeMux I__674 (
            .O(N__4231),
            .I(N__4220));
    CascadeMux I__673 (
            .O(N__4230),
            .I(N__4217));
    Span4Mux_s3_h I__672 (
            .O(N__4227),
            .I(N__4214));
    LocalMux I__671 (
            .O(N__4224),
            .I(N__4211));
    InMux I__670 (
            .O(N__4223),
            .I(N__4204));
    InMux I__669 (
            .O(N__4220),
            .I(N__4204));
    InMux I__668 (
            .O(N__4217),
            .I(N__4204));
    Odrv4 I__667 (
            .O(N__4214),
            .I(r_CountZ0Z_3));
    Odrv4 I__666 (
            .O(N__4211),
            .I(r_CountZ0Z_3));
    LocalMux I__665 (
            .O(N__4204),
            .I(r_CountZ0Z_3));
    InMux I__664 (
            .O(N__4197),
            .I(N__4194));
    LocalMux I__663 (
            .O(N__4194),
            .I(N__4191));
    Odrv4 I__662 (
            .O(N__4191),
            .I(sevsegl_RNO_0Z0Z_3));
    InMux I__661 (
            .O(N__4188),
            .I(N__4184));
    CascadeMux I__660 (
            .O(N__4187),
            .I(N__4179));
    LocalMux I__659 (
            .O(N__4184),
            .I(N__4174));
    InMux I__658 (
            .O(N__4183),
            .I(N__4171));
    InMux I__657 (
            .O(N__4182),
            .I(N__4164));
    InMux I__656 (
            .O(N__4179),
            .I(N__4164));
    InMux I__655 (
            .O(N__4178),
            .I(N__4164));
    CascadeMux I__654 (
            .O(N__4177),
            .I(N__4161));
    Span4Mux_s3_h I__653 (
            .O(N__4174),
            .I(N__4157));
    LocalMux I__652 (
            .O(N__4171),
            .I(N__4154));
    LocalMux I__651 (
            .O(N__4164),
            .I(N__4151));
    InMux I__650 (
            .O(N__4161),
            .I(N__4146));
    InMux I__649 (
            .O(N__4160),
            .I(N__4146));
    Odrv4 I__648 (
            .O(N__4157),
            .I(\alogicunit.result24 ));
    Odrv4 I__647 (
            .O(N__4154),
            .I(\alogicunit.result24 ));
    Odrv4 I__646 (
            .O(N__4151),
            .I(\alogicunit.result24 ));
    LocalMux I__645 (
            .O(N__4146),
            .I(\alogicunit.result24 ));
    CascadeMux I__644 (
            .O(N__4137),
            .I(\alogicunit.result24_cascade_ ));
    CascadeMux I__643 (
            .O(N__4134),
            .I(N__4130));
    InMux I__642 (
            .O(N__4133),
            .I(N__4126));
    InMux I__641 (
            .O(N__4130),
            .I(N__4123));
    InMux I__640 (
            .O(N__4129),
            .I(N__4120));
    LocalMux I__639 (
            .O(N__4126),
            .I(N__4117));
    LocalMux I__638 (
            .O(N__4123),
            .I(N__4114));
    LocalMux I__637 (
            .O(N__4120),
            .I(\alogicunit.un1_a_1_axb_3 ));
    Odrv4 I__636 (
            .O(N__4117),
            .I(\alogicunit.un1_a_1_axb_3 ));
    Odrv4 I__635 (
            .O(N__4114),
            .I(\alogicunit.un1_a_1_axb_3 ));
    CascadeMux I__634 (
            .O(N__4107),
            .I(N__4103));
    CascadeMux I__633 (
            .O(N__4106),
            .I(N__4100));
    InMux I__632 (
            .O(N__4103),
            .I(N__4095));
    InMux I__631 (
            .O(N__4100),
            .I(N__4095));
    LocalMux I__630 (
            .O(N__4095),
            .I(N__4092));
    Span12Mux_s3_h I__629 (
            .O(N__4092),
            .I(N__4089));
    Odrv12 I__628 (
            .O(N__4089),
            .I(\alogicunit.N_51 ));
    InMux I__627 (
            .O(N__4086),
            .I(N__4080));
    InMux I__626 (
            .O(N__4085),
            .I(N__4080));
    LocalMux I__625 (
            .O(N__4080),
            .I(cu1_track_ns_3));
    CascadeMux I__624 (
            .O(N__4077),
            .I(N__4074));
    InMux I__623 (
            .O(N__4074),
            .I(N__4071));
    LocalMux I__622 (
            .O(N__4071),
            .I(\alogicunit.un1_a_1_cry_1_THRU_CO ));
    InMux I__621 (
            .O(N__4068),
            .I(\alogicunit.un1_a_1_cry_1 ));
    InMux I__620 (
            .O(N__4065),
            .I(N__4062));
    LocalMux I__619 (
            .O(N__4062),
            .I(\alogicunit.un1_a_1_cry_2_THRU_CO ));
    InMux I__618 (
            .O(N__4059),
            .I(\alogicunit.un1_a_1_cry_2 ));
    InMux I__617 (
            .O(N__4056),
            .I(\alogicunit.un1_a_1_cry_3 ));
    InMux I__616 (
            .O(N__4053),
            .I(N__4050));
    LocalMux I__615 (
            .O(N__4050),
            .I(N__4047));
    Odrv4 I__614 (
            .O(N__4047),
            .I(\alogicunit.result_RNO_0Z0Z_5 ));
    InMux I__613 (
            .O(N__4044),
            .I(\alogicunit.un1_a_1_cry_4 ));
    InMux I__612 (
            .O(N__4041),
            .I(\alogicunit.un1_a_1_cry_5 ));
    CascadeMux I__611 (
            .O(N__4038),
            .I(N__4033));
    InMux I__610 (
            .O(N__4037),
            .I(N__4028));
    InMux I__609 (
            .O(N__4036),
            .I(N__4028));
    InMux I__608 (
            .O(N__4033),
            .I(N__4025));
    LocalMux I__607 (
            .O(N__4028),
            .I(\alogicunit.N_95_1 ));
    LocalMux I__606 (
            .O(N__4025),
            .I(\alogicunit.N_95_1 ));
    InMux I__605 (
            .O(N__4020),
            .I(\alogicunit.un1_a_1_cry_6 ));
    InMux I__604 (
            .O(N__4017),
            .I(N__4014));
    LocalMux I__603 (
            .O(N__4014),
            .I(N__4011));
    Odrv4 I__602 (
            .O(N__4011),
            .I(left_3));
    CascadeMux I__601 (
            .O(N__4008),
            .I(N__4005));
    InMux I__600 (
            .O(N__4005),
            .I(N__4002));
    LocalMux I__599 (
            .O(N__4002),
            .I(\alogicunit.m26_l_fxZ0Z_0 ));
    CascadeMux I__598 (
            .O(N__3999),
            .I(un1_click13_1_sn_cascade_));
    InMux I__597 (
            .O(N__3996),
            .I(N__3993));
    LocalMux I__596 (
            .O(N__3993),
            .I(N__3990));
    Odrv12 I__595 (
            .O(N__3990),
            .I(sevsegr_RNO_0Z0Z_2));
    InMux I__594 (
            .O(N__3987),
            .I(N__3984));
    LocalMux I__593 (
            .O(N__3984),
            .I(N__3979));
    InMux I__592 (
            .O(N__3983),
            .I(N__3976));
    InMux I__591 (
            .O(N__3982),
            .I(N__3973));
    Span4Mux_s3_h I__590 (
            .O(N__3979),
            .I(N__3970));
    LocalMux I__589 (
            .O(N__3976),
            .I(r_Count11));
    LocalMux I__588 (
            .O(N__3973),
            .I(r_Count11));
    Odrv4 I__587 (
            .O(N__3970),
            .I(r_Count11));
    CascadeMux I__586 (
            .O(N__3963),
            .I(r_Count11_cascade_));
    CascadeMux I__585 (
            .O(N__3960),
            .I(\alogicunit.N_95_1_cascade_ ));
    CascadeMux I__584 (
            .O(N__3957),
            .I(N__3954));
    InMux I__583 (
            .O(N__3954),
            .I(N__3951));
    LocalMux I__582 (
            .O(N__3951),
            .I(N__3948));
    Span4Mux_s3_h I__581 (
            .O(N__3948),
            .I(N__3945));
    Odrv4 I__580 (
            .O(N__3945),
            .I(right_0));
    InMux I__579 (
            .O(N__3942),
            .I(N__3939));
    LocalMux I__578 (
            .O(N__3939),
            .I(right_3));
    InMux I__577 (
            .O(N__3936),
            .I(N__3933));
    LocalMux I__576 (
            .O(N__3933),
            .I(N__3930));
    Span4Mux_s3_h I__575 (
            .O(N__3930),
            .I(N__3926));
    InMux I__574 (
            .O(N__3929),
            .I(N__3923));
    Odrv4 I__573 (
            .O(N__3926),
            .I(SUM_3));
    LocalMux I__572 (
            .O(N__3923),
            .I(SUM_3));
    InMux I__571 (
            .O(N__3918),
            .I(N__3915));
    LocalMux I__570 (
            .O(N__3915),
            .I(N__3912));
    Span4Mux_v I__569 (
            .O(N__3912),
            .I(N__3909));
    Odrv4 I__568 (
            .O(N__3909),
            .I(sevsegr_RNO_1Z0Z_3));
    InMux I__567 (
            .O(N__3906),
            .I(N__3903));
    LocalMux I__566 (
            .O(N__3903),
            .I(N__3900));
    Span4Mux_s3_h I__565 (
            .O(N__3900),
            .I(N__3897));
    Odrv4 I__564 (
            .O(N__3897),
            .I(right_2));
    InMux I__563 (
            .O(N__3894),
            .I(N__3891));
    LocalMux I__562 (
            .O(N__3891),
            .I(sevsegl_7_ns_1_0));
    InMux I__561 (
            .O(N__3888),
            .I(N__3864));
    InMux I__560 (
            .O(N__3887),
            .I(N__3864));
    InMux I__559 (
            .O(N__3886),
            .I(N__3864));
    InMux I__558 (
            .O(N__3885),
            .I(N__3864));
    InMux I__557 (
            .O(N__3884),
            .I(N__3864));
    InMux I__556 (
            .O(N__3883),
            .I(N__3864));
    InMux I__555 (
            .O(N__3882),
            .I(N__3864));
    InMux I__554 (
            .O(N__3881),
            .I(N__3861));
    InMux I__553 (
            .O(N__3880),
            .I(N__3858));
    InMux I__552 (
            .O(N__3879),
            .I(N__3855));
    LocalMux I__551 (
            .O(N__3864),
            .I(r_Switch_2_RNIK7AZ0Z11));
    LocalMux I__550 (
            .O(N__3861),
            .I(r_Switch_2_RNIK7AZ0Z11));
    LocalMux I__549 (
            .O(N__3858),
            .I(r_Switch_2_RNIK7AZ0Z11));
    LocalMux I__548 (
            .O(N__3855),
            .I(r_Switch_2_RNIK7AZ0Z11));
    CEMux I__547 (
            .O(N__3846),
            .I(N__3843));
    LocalMux I__546 (
            .O(N__3843),
            .I(N__3839));
    CEMux I__545 (
            .O(N__3842),
            .I(N__3836));
    Span4Mux_h I__544 (
            .O(N__3839),
            .I(N__3833));
    LocalMux I__543 (
            .O(N__3836),
            .I(N__3830));
    Odrv4 I__542 (
            .O(N__3833),
            .I(un1_click17_0));
    Odrv4 I__541 (
            .O(N__3830),
            .I(un1_click17_0));
    IoInMux I__540 (
            .O(N__3825),
            .I(N__3822));
    LocalMux I__539 (
            .O(N__3822),
            .I(r_HexEncode_i_4));
    IoInMux I__538 (
            .O(N__3819),
            .I(N__3816));
    LocalMux I__537 (
            .O(N__3816),
            .I(N__3813));
    IoSpan4Mux I__536 (
            .O(N__3813),
            .I(N__3810));
    Span4Mux_s0_v I__535 (
            .O(N__3810),
            .I(N__3807));
    Odrv4 I__534 (
            .O(N__3807),
            .I(r_HexEncode_i_0));
    IoInMux I__533 (
            .O(N__3804),
            .I(N__3801));
    LocalMux I__532 (
            .O(N__3801),
            .I(N__3798));
    IoSpan4Mux I__531 (
            .O(N__3798),
            .I(N__3795));
    Odrv4 I__530 (
            .O(N__3795),
            .I(r_HexEncode_i_2));
    IoInMux I__529 (
            .O(N__3792),
            .I(N__3789));
    LocalMux I__528 (
            .O(N__3789),
            .I(N__3786));
    IoSpan4Mux I__527 (
            .O(N__3786),
            .I(N__3783));
    Odrv4 I__526 (
            .O(N__3783),
            .I(r_HexEncode_i_3));
    CascadeMux I__525 (
            .O(N__3780),
            .I(N__3777));
    InMux I__524 (
            .O(N__3777),
            .I(N__3774));
    LocalMux I__523 (
            .O(N__3774),
            .I(N__3765));
    InMux I__522 (
            .O(N__3773),
            .I(N__3754));
    InMux I__521 (
            .O(N__3772),
            .I(N__3754));
    InMux I__520 (
            .O(N__3771),
            .I(N__3754));
    InMux I__519 (
            .O(N__3770),
            .I(N__3754));
    InMux I__518 (
            .O(N__3769),
            .I(N__3754));
    InMux I__517 (
            .O(N__3768),
            .I(N__3751));
    Span4Mux_s1_h I__516 (
            .O(N__3765),
            .I(N__3746));
    LocalMux I__515 (
            .O(N__3754),
            .I(N__3746));
    LocalMux I__514 (
            .O(N__3751),
            .I(sevsegrZ0Z_0));
    Odrv4 I__513 (
            .O(N__3746),
            .I(sevsegrZ0Z_0));
    InMux I__512 (
            .O(N__3741),
            .I(N__3733));
    InMux I__511 (
            .O(N__3740),
            .I(N__3722));
    InMux I__510 (
            .O(N__3739),
            .I(N__3722));
    InMux I__509 (
            .O(N__3738),
            .I(N__3722));
    InMux I__508 (
            .O(N__3737),
            .I(N__3722));
    InMux I__507 (
            .O(N__3736),
            .I(N__3722));
    LocalMux I__506 (
            .O(N__3733),
            .I(N__3716));
    LocalMux I__505 (
            .O(N__3722),
            .I(N__3716));
    InMux I__504 (
            .O(N__3721),
            .I(N__3713));
    Odrv4 I__503 (
            .O(N__3716),
            .I(sevsegrZ0Z_2));
    LocalMux I__502 (
            .O(N__3713),
            .I(sevsegrZ0Z_2));
    InMux I__501 (
            .O(N__3708),
            .I(N__3702));
    CascadeMux I__500 (
            .O(N__3707),
            .I(N__3699));
    CascadeMux I__499 (
            .O(N__3706),
            .I(N__3696));
    CascadeMux I__498 (
            .O(N__3705),
            .I(N__3692));
    LocalMux I__497 (
            .O(N__3702),
            .I(N__3688));
    InMux I__496 (
            .O(N__3699),
            .I(N__3677));
    InMux I__495 (
            .O(N__3696),
            .I(N__3677));
    InMux I__494 (
            .O(N__3695),
            .I(N__3677));
    InMux I__493 (
            .O(N__3692),
            .I(N__3677));
    InMux I__492 (
            .O(N__3691),
            .I(N__3677));
    Sp12to4 I__491 (
            .O(N__3688),
            .I(N__3671));
    LocalMux I__490 (
            .O(N__3677),
            .I(N__3671));
    InMux I__489 (
            .O(N__3676),
            .I(N__3668));
    Odrv12 I__488 (
            .O(N__3671),
            .I(sevsegrZ0Z_1));
    LocalMux I__487 (
            .O(N__3668),
            .I(sevsegrZ0Z_1));
    CascadeMux I__486 (
            .O(N__3663),
            .I(N__3656));
    CascadeMux I__485 (
            .O(N__3662),
            .I(N__3652));
    InMux I__484 (
            .O(N__3661),
            .I(N__3648));
    InMux I__483 (
            .O(N__3660),
            .I(N__3637));
    InMux I__482 (
            .O(N__3659),
            .I(N__3637));
    InMux I__481 (
            .O(N__3656),
            .I(N__3637));
    InMux I__480 (
            .O(N__3655),
            .I(N__3637));
    InMux I__479 (
            .O(N__3652),
            .I(N__3637));
    CascadeMux I__478 (
            .O(N__3651),
            .I(N__3634));
    LocalMux I__477 (
            .O(N__3648),
            .I(N__3629));
    LocalMux I__476 (
            .O(N__3637),
            .I(N__3629));
    InMux I__475 (
            .O(N__3634),
            .I(N__3626));
    Odrv4 I__474 (
            .O(N__3629),
            .I(sevsegrZ0Z_3));
    LocalMux I__473 (
            .O(N__3626),
            .I(sevsegrZ0Z_3));
    IoInMux I__472 (
            .O(N__3621),
            .I(N__3618));
    LocalMux I__471 (
            .O(N__3618),
            .I(r_HexEncode_i_5));
    CascadeMux I__470 (
            .O(N__3615),
            .I(SUM_3_cascade_));
    InMux I__469 (
            .O(N__3612),
            .I(N__3609));
    LocalMux I__468 (
            .O(N__3609),
            .I(sevsegl_RNO_1Z0Z_3));
    InMux I__467 (
            .O(N__3606),
            .I(N__3603));
    LocalMux I__466 (
            .O(N__3603),
            .I(N__3600));
    Odrv4 I__465 (
            .O(N__3600),
            .I(sevsegr_RNO_1Z0Z_1));
    CascadeMux I__464 (
            .O(N__3597),
            .I(N__3594));
    InMux I__463 (
            .O(N__3594),
            .I(N__3591));
    LocalMux I__462 (
            .O(N__3591),
            .I(sevsegr_RNO_1Z0Z_2));
    InMux I__461 (
            .O(N__3588),
            .I(N__3585));
    LocalMux I__460 (
            .O(N__3585),
            .I(N__3582));
    Odrv4 I__459 (
            .O(N__3582),
            .I(sevsegr_RNO_0Z0Z_3));
    InMux I__458 (
            .O(N__3579),
            .I(N__3576));
    LocalMux I__457 (
            .O(N__3576),
            .I(sevsegl_RNO_1Z0Z_1));
    InMux I__456 (
            .O(N__3573),
            .I(N__3570));
    LocalMux I__455 (
            .O(N__3570),
            .I(sevsegr_7_ns_1_0));
    CascadeMux I__454 (
            .O(N__3567),
            .I(N__3562));
    InMux I__453 (
            .O(N__3566),
            .I(N__3559));
    InMux I__452 (
            .O(N__3565),
            .I(N__3556));
    InMux I__451 (
            .O(N__3562),
            .I(N__3553));
    LocalMux I__450 (
            .O(N__3559),
            .I(\Instance1.r_CountZ0Z_14 ));
    LocalMux I__449 (
            .O(N__3556),
            .I(\Instance1.r_CountZ0Z_14 ));
    LocalMux I__448 (
            .O(N__3553),
            .I(\Instance1.r_CountZ0Z_14 ));
    InMux I__447 (
            .O(N__3546),
            .I(\Instance1.r_Count_2_cry_13 ));
    InMux I__446 (
            .O(N__3543),
            .I(N__3538));
    InMux I__445 (
            .O(N__3542),
            .I(N__3535));
    InMux I__444 (
            .O(N__3541),
            .I(N__3532));
    LocalMux I__443 (
            .O(N__3538),
            .I(\Instance1.r_CountZ0Z_15 ));
    LocalMux I__442 (
            .O(N__3535),
            .I(\Instance1.r_CountZ0Z_15 ));
    LocalMux I__441 (
            .O(N__3532),
            .I(\Instance1.r_CountZ0Z_15 ));
    InMux I__440 (
            .O(N__3525),
            .I(\Instance1.r_Count_2_cry_14 ));
    CascadeMux I__439 (
            .O(N__3522),
            .I(N__3518));
    InMux I__438 (
            .O(N__3521),
            .I(N__3514));
    InMux I__437 (
            .O(N__3518),
            .I(N__3511));
    InMux I__436 (
            .O(N__3517),
            .I(N__3508));
    LocalMux I__435 (
            .O(N__3514),
            .I(\Instance1.r_CountZ0Z_16 ));
    LocalMux I__434 (
            .O(N__3511),
            .I(\Instance1.r_CountZ0Z_16 ));
    LocalMux I__433 (
            .O(N__3508),
            .I(\Instance1.r_CountZ0Z_16 ));
    InMux I__432 (
            .O(N__3501),
            .I(\Instance1.r_Count_2_cry_15 ));
    InMux I__431 (
            .O(N__3498),
            .I(bfn_2_11_0_));
    InMux I__430 (
            .O(N__3495),
            .I(N__3490));
    InMux I__429 (
            .O(N__3494),
            .I(N__3487));
    InMux I__428 (
            .O(N__3493),
            .I(N__3484));
    LocalMux I__427 (
            .O(N__3490),
            .I(\Instance1.r_CountZ0Z_17 ));
    LocalMux I__426 (
            .O(N__3487),
            .I(\Instance1.r_CountZ0Z_17 ));
    LocalMux I__425 (
            .O(N__3484),
            .I(\Instance1.r_CountZ0Z_17 ));
    CascadeMux I__424 (
            .O(N__3477),
            .I(N__3474));
    InMux I__423 (
            .O(N__3474),
            .I(N__3468));
    InMux I__422 (
            .O(N__3473),
            .I(N__3465));
    InMux I__421 (
            .O(N__3472),
            .I(N__3462));
    InMux I__420 (
            .O(N__3471),
            .I(N__3459));
    LocalMux I__419 (
            .O(N__3468),
            .I(N__3456));
    LocalMux I__418 (
            .O(N__3465),
            .I(\Instance1.r_CountZ0Z_0 ));
    LocalMux I__417 (
            .O(N__3462),
            .I(\Instance1.r_CountZ0Z_0 ));
    LocalMux I__416 (
            .O(N__3459),
            .I(\Instance1.r_CountZ0Z_0 ));
    Odrv4 I__415 (
            .O(N__3456),
            .I(\Instance1.r_CountZ0Z_0 ));
    SRMux I__414 (
            .O(N__3447),
            .I(N__3435));
    SRMux I__413 (
            .O(N__3446),
            .I(N__3435));
    SRMux I__412 (
            .O(N__3445),
            .I(N__3435));
    SRMux I__411 (
            .O(N__3444),
            .I(N__3435));
    GlobalMux I__410 (
            .O(N__3435),
            .I(N__3432));
    gio2CtrlBuf I__409 (
            .O(N__3432),
            .I(\Instance1.r_Count12_i_g ));
    CascadeMux I__408 (
            .O(N__3429),
            .I(N__3426));
    InMux I__407 (
            .O(N__3426),
            .I(N__3423));
    LocalMux I__406 (
            .O(N__3423),
            .I(left_1));
    CascadeMux I__405 (
            .O(N__3420),
            .I(N__3417));
    InMux I__404 (
            .O(N__3417),
            .I(N__3414));
    LocalMux I__403 (
            .O(N__3414),
            .I(right_1));
    InMux I__402 (
            .O(N__3411),
            .I(N__3406));
    InMux I__401 (
            .O(N__3410),
            .I(N__3401));
    InMux I__400 (
            .O(N__3409),
            .I(N__3401));
    LocalMux I__399 (
            .O(N__3406),
            .I(\Instance1.r_CountZ0Z_6 ));
    LocalMux I__398 (
            .O(N__3401),
            .I(\Instance1.r_CountZ0Z_6 ));
    InMux I__397 (
            .O(N__3396),
            .I(\Instance1.r_Count_2_cry_5 ));
    CascadeMux I__396 (
            .O(N__3393),
            .I(N__3388));
    InMux I__395 (
            .O(N__3392),
            .I(N__3385));
    InMux I__394 (
            .O(N__3391),
            .I(N__3380));
    InMux I__393 (
            .O(N__3388),
            .I(N__3380));
    LocalMux I__392 (
            .O(N__3385),
            .I(N__3375));
    LocalMux I__391 (
            .O(N__3380),
            .I(N__3375));
    Odrv4 I__390 (
            .O(N__3375),
            .I(\Instance1.r_CountZ0Z_7 ));
    InMux I__389 (
            .O(N__3372),
            .I(\Instance1.r_Count_2_cry_6 ));
    InMux I__388 (
            .O(N__3369),
            .I(N__3364));
    InMux I__387 (
            .O(N__3368),
            .I(N__3359));
    InMux I__386 (
            .O(N__3367),
            .I(N__3359));
    LocalMux I__385 (
            .O(N__3364),
            .I(\Instance1.r_CountZ0Z_8 ));
    LocalMux I__384 (
            .O(N__3359),
            .I(\Instance1.r_CountZ0Z_8 ));
    InMux I__383 (
            .O(N__3354),
            .I(\Instance1.r_Count_2_cry_7 ));
    CascadeMux I__382 (
            .O(N__3351),
            .I(N__3346));
    InMux I__381 (
            .O(N__3350),
            .I(N__3343));
    InMux I__380 (
            .O(N__3349),
            .I(N__3340));
    InMux I__379 (
            .O(N__3346),
            .I(N__3337));
    LocalMux I__378 (
            .O(N__3343),
            .I(\Instance1.r_CountZ0Z_9 ));
    LocalMux I__377 (
            .O(N__3340),
            .I(\Instance1.r_CountZ0Z_9 ));
    LocalMux I__376 (
            .O(N__3337),
            .I(\Instance1.r_CountZ0Z_9 ));
    InMux I__375 (
            .O(N__3330),
            .I(bfn_2_10_0_));
    CascadeMux I__374 (
            .O(N__3327),
            .I(N__3324));
    InMux I__373 (
            .O(N__3324),
            .I(N__3319));
    InMux I__372 (
            .O(N__3323),
            .I(N__3316));
    InMux I__371 (
            .O(N__3322),
            .I(N__3313));
    LocalMux I__370 (
            .O(N__3319),
            .I(\Instance1.r_CountZ0Z_10 ));
    LocalMux I__369 (
            .O(N__3316),
            .I(\Instance1.r_CountZ0Z_10 ));
    LocalMux I__368 (
            .O(N__3313),
            .I(\Instance1.r_CountZ0Z_10 ));
    InMux I__367 (
            .O(N__3306),
            .I(\Instance1.r_Count_2_cry_9 ));
    InMux I__366 (
            .O(N__3303),
            .I(N__3298));
    InMux I__365 (
            .O(N__3302),
            .I(N__3295));
    InMux I__364 (
            .O(N__3301),
            .I(N__3292));
    LocalMux I__363 (
            .O(N__3298),
            .I(\Instance1.r_CountZ0Z_11 ));
    LocalMux I__362 (
            .O(N__3295),
            .I(\Instance1.r_CountZ0Z_11 ));
    LocalMux I__361 (
            .O(N__3292),
            .I(\Instance1.r_CountZ0Z_11 ));
    InMux I__360 (
            .O(N__3285),
            .I(\Instance1.r_Count_2_cry_10 ));
    CascadeMux I__359 (
            .O(N__3282),
            .I(N__3278));
    InMux I__358 (
            .O(N__3281),
            .I(N__3274));
    InMux I__357 (
            .O(N__3278),
            .I(N__3269));
    InMux I__356 (
            .O(N__3277),
            .I(N__3269));
    LocalMux I__355 (
            .O(N__3274),
            .I(\Instance1.r_CountZ0Z_12 ));
    LocalMux I__354 (
            .O(N__3269),
            .I(\Instance1.r_CountZ0Z_12 ));
    InMux I__353 (
            .O(N__3264),
            .I(\Instance1.r_Count_2_cry_11 ));
    InMux I__352 (
            .O(N__3261),
            .I(N__3256));
    InMux I__351 (
            .O(N__3260),
            .I(N__3251));
    InMux I__350 (
            .O(N__3259),
            .I(N__3251));
    LocalMux I__349 (
            .O(N__3256),
            .I(\Instance1.r_CountZ0Z_13 ));
    LocalMux I__348 (
            .O(N__3251),
            .I(\Instance1.r_CountZ0Z_13 ));
    InMux I__347 (
            .O(N__3246),
            .I(\Instance1.r_Count_2_cry_12 ));
    CascadeMux I__346 (
            .O(N__3243),
            .I(SUM_2_cascade_));
    IoInMux I__345 (
            .O(N__3240),
            .I(N__3237));
    LocalMux I__344 (
            .O(N__3237),
            .I(r_HexEncode_i_0_0));
    IoInMux I__343 (
            .O(N__3234),
            .I(N__3231));
    LocalMux I__342 (
            .O(N__3231),
            .I(r_HexEncode_i_0_1));
    IoInMux I__341 (
            .O(N__3228),
            .I(N__3225));
    LocalMux I__340 (
            .O(N__3225),
            .I(r_HexEncode_i_6));
    InMux I__339 (
            .O(N__3222),
            .I(N__3217));
    InMux I__338 (
            .O(N__3221),
            .I(N__3212));
    InMux I__337 (
            .O(N__3220),
            .I(N__3212));
    LocalMux I__336 (
            .O(N__3217),
            .I(\Instance1.r_CountZ0Z_1 ));
    LocalMux I__335 (
            .O(N__3212),
            .I(\Instance1.r_CountZ0Z_1 ));
    InMux I__334 (
            .O(N__3207),
            .I(N__3203));
    InMux I__333 (
            .O(N__3206),
            .I(N__3200));
    LocalMux I__332 (
            .O(N__3203),
            .I(\Instance1.r_CountZ0Z_2 ));
    LocalMux I__331 (
            .O(N__3200),
            .I(\Instance1.r_CountZ0Z_2 ));
    InMux I__330 (
            .O(N__3195),
            .I(\Instance1.r_Count_2_cry_1 ));
    CascadeMux I__329 (
            .O(N__3192),
            .I(N__3188));
    InMux I__328 (
            .O(N__3191),
            .I(N__3185));
    InMux I__327 (
            .O(N__3188),
            .I(N__3182));
    LocalMux I__326 (
            .O(N__3185),
            .I(\Instance1.r_CountZ0Z_3 ));
    LocalMux I__325 (
            .O(N__3182),
            .I(\Instance1.r_CountZ0Z_3 ));
    InMux I__324 (
            .O(N__3177),
            .I(\Instance1.r_Count_2_cry_2 ));
    InMux I__323 (
            .O(N__3174),
            .I(N__3169));
    InMux I__322 (
            .O(N__3173),
            .I(N__3166));
    InMux I__321 (
            .O(N__3172),
            .I(N__3163));
    LocalMux I__320 (
            .O(N__3169),
            .I(N__3158));
    LocalMux I__319 (
            .O(N__3166),
            .I(N__3158));
    LocalMux I__318 (
            .O(N__3163),
            .I(\Instance1.r_CountZ0Z_4 ));
    Odrv12 I__317 (
            .O(N__3158),
            .I(\Instance1.r_CountZ0Z_4 ));
    InMux I__316 (
            .O(N__3153),
            .I(\Instance1.r_Count_2_cry_3 ));
    InMux I__315 (
            .O(N__3150),
            .I(N__3147));
    LocalMux I__314 (
            .O(N__3147),
            .I(N__3142));
    InMux I__313 (
            .O(N__3146),
            .I(N__3139));
    InMux I__312 (
            .O(N__3145),
            .I(N__3136));
    Odrv4 I__311 (
            .O(N__3142),
            .I(\Instance1.r_CountZ0Z_5 ));
    LocalMux I__310 (
            .O(N__3139),
            .I(\Instance1.r_CountZ0Z_5 ));
    LocalMux I__309 (
            .O(N__3136),
            .I(\Instance1.r_CountZ0Z_5 ));
    InMux I__308 (
            .O(N__3129),
            .I(\Instance1.r_Count_2_cry_4 ));
    CascadeMux I__307 (
            .O(N__3126),
            .I(sevsegl_RNO_0Z0Z_2_cascade_));
    InMux I__306 (
            .O(N__3123),
            .I(N__3120));
    LocalMux I__305 (
            .O(N__3120),
            .I(sevsegl_RNO_1Z0Z_2));
    IoInMux I__304 (
            .O(N__3117),
            .I(N__3114));
    LocalMux I__303 (
            .O(N__3114),
            .I(r_HexEncode_i_0_6));
    IoInMux I__302 (
            .O(N__3111),
            .I(N__3108));
    LocalMux I__301 (
            .O(N__3108),
            .I(r_HexEncode_i_1));
    IoInMux I__300 (
            .O(N__3105),
            .I(N__3102));
    LocalMux I__299 (
            .O(N__3102),
            .I(r_HexEncode_i_0_5));
    InMux I__298 (
            .O(N__3099),
            .I(N__3096));
    LocalMux I__297 (
            .O(N__3096),
            .I(SUM_2));
    InMux I__296 (
            .O(N__3093),
            .I(N__3090));
    LocalMux I__295 (
            .O(N__3090),
            .I(\Instance1.un1_r_Count_10lto17_1 ));
    InMux I__294 (
            .O(N__3087),
            .I(N__3084));
    LocalMux I__293 (
            .O(N__3084),
            .I(r_SwitchZ0Z_1));
    InMux I__292 (
            .O(N__3081),
            .I(N__3078));
    LocalMux I__291 (
            .O(N__3078),
            .I(N__3075));
    Odrv4 I__290 (
            .O(N__3075),
            .I(\Instance1.r_Count13_8_0 ));
    CascadeMux I__289 (
            .O(N__3072),
            .I(\Instance1.r_Count13_4_cascade_ ));
    InMux I__288 (
            .O(N__3069),
            .I(N__3066));
    LocalMux I__287 (
            .O(N__3066),
            .I(\Instance1.r_Count13_7 ));
    InMux I__286 (
            .O(N__3063),
            .I(N__3060));
    LocalMux I__285 (
            .O(N__3060),
            .I(N__3057));
    Odrv4 I__284 (
            .O(N__3057),
            .I(\Instance1.r_Count13_10 ));
    InMux I__283 (
            .O(N__3054),
            .I(N__3050));
    InMux I__282 (
            .O(N__3053),
            .I(N__3047));
    LocalMux I__281 (
            .O(N__3050),
            .I(N__3044));
    LocalMux I__280 (
            .O(N__3047),
            .I(N__3041));
    Span4Mux_v I__279 (
            .O(N__3044),
            .I(N__3038));
    Sp12to4 I__278 (
            .O(N__3041),
            .I(N__3033));
    Sp12to4 I__277 (
            .O(N__3038),
            .I(N__3033));
    Span12Mux_v I__276 (
            .O(N__3033),
            .I(N__3030));
    Odrv12 I__275 (
            .O(N__3030),
            .I(i_Switch_1_c));
    InMux I__274 (
            .O(N__3027),
            .I(N__3024));
    LocalMux I__273 (
            .O(N__3024),
            .I(\Instance1.r_Count13_12 ));
    CascadeMux I__272 (
            .O(N__3021),
            .I(\Instance1.r_Count13_13_cascade_ ));
    InMux I__271 (
            .O(N__3018),
            .I(N__3015));
    LocalMux I__270 (
            .O(N__3015),
            .I(N__3009));
    InMux I__269 (
            .O(N__3014),
            .I(N__3002));
    InMux I__268 (
            .O(N__3013),
            .I(N__3002));
    InMux I__267 (
            .O(N__3012),
            .I(N__3002));
    Odrv12 I__266 (
            .O(N__3009),
            .I(w_Switch_1));
    LocalMux I__265 (
            .O(N__3002),
            .I(w_Switch_1));
    CascadeMux I__264 (
            .O(N__2997),
            .I(\Instance1.un1_r_Count_10lt11_0_cascade_ ));
    InMux I__263 (
            .O(N__2994),
            .I(N__2991));
    LocalMux I__262 (
            .O(N__2991),
            .I(\Instance1.un1_r_Count_10lto11_1 ));
    CascadeMux I__261 (
            .O(N__2988),
            .I(\Instance1.un1_r_Count_10lt17_cascade_ ));
    IoInMux I__260 (
            .O(N__2985),
            .I(N__2982));
    LocalMux I__259 (
            .O(N__2982),
            .I(\Instance1.r_Count12_i ));
    defparam IN_MUX_bfv_4_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_12_0_));
    defparam IN_MUX_bfv_6_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_7_0_));
    defparam IN_MUX_bfv_6_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_8_0_ (
            .carryinitin(\Instance4.r_Count_2_cry_8 ),
            .carryinitout(bfn_6_8_0_));
    defparam IN_MUX_bfv_6_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_9_0_ (
            .carryinitin(\Instance4.r_Count_2_cry_16 ),
            .carryinitout(bfn_6_9_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(\Instance3.r_Count_2_cry_8 ),
            .carryinitout(bfn_8_10_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(\Instance3.r_Count_2_cry_16 ),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_6_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_10_0_));
    defparam IN_MUX_bfv_6_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_11_0_ (
            .carryinitin(\Instance2.r_Count_2_cry_8 ),
            .carryinitout(bfn_6_11_0_));
    defparam IN_MUX_bfv_6_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_12_0_ (
            .carryinitin(\Instance2.r_Count_2_cry_16 ),
            .carryinitout(bfn_6_12_0_));
    defparam IN_MUX_bfv_2_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_9_0_));
    defparam IN_MUX_bfv_2_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_10_0_ (
            .carryinitin(\Instance1.r_Count_2_cry_8 ),
            .carryinitout(bfn_2_10_0_));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(\Instance1.r_Count_2_cry_16 ),
            .carryinitout(bfn_2_11_0_));
    ICE_GB \Instance1.r_State_RNIK9757_0  (
            .USERSIGNALTOGLOBALBUFFER(N__2985),
            .GLOBALBUFFEROUTPUT(\Instance1.r_Count12_i_g ));
    ICE_GB \Instance4.r_State_RNI4ONP3_0  (
            .USERSIGNALTOGLOBALBUFFER(N__6204),
            .GLOBALBUFFEROUTPUT(\Instance4.r_Count12_i_g ));
    ICE_GB \Instance2.r_State_RNI4PC15_0  (
            .USERSIGNALTOGLOBALBUFFER(N__4839),
            .GLOBALBUFFEROUTPUT(\Instance2.r_Count12_i_g ));
    ICE_GB \Instance3.r_State_RNIK8IT5_0  (
            .USERSIGNALTOGLOBALBUFFER(N__6498),
            .GLOBALBUFFEROUTPUT(\Instance3.r_Count12_i_g ));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \Instance1.r_State_RNO_5_LC_1_9_1 .C_ON=1'b0;
    defparam \Instance1.r_State_RNO_5_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \Instance1.r_State_RNO_5_LC_1_9_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Instance1.r_State_RNO_5_LC_1_9_1  (
            .in0(N__3410),
            .in1(N__3542),
            .in2(N__3522),
            .in3(N__3368),
            .lcout(\Instance1.r_Count13_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance1.r_Count_RNIC2TU1_8_LC_1_9_3 .C_ON=1'b0;
    defparam \Instance1.r_Count_RNIC2TU1_8_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \Instance1.r_Count_RNIC2TU1_8_LC_1_9_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Instance1.r_Count_RNIC2TU1_8_LC_1_9_3  (
            .in0(N__3322),
            .in1(N__3301),
            .in2(N__3351),
            .in3(N__3367),
            .lcout(\Instance1.un1_r_Count_10lto11_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance1.r_Count_RNIED2U1_4_LC_1_9_4 .C_ON=1'b0;
    defparam \Instance1.r_Count_RNIED2U1_4_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \Instance1.r_Count_RNIED2U1_4_LC_1_9_4 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \Instance1.r_Count_RNIED2U1_4_LC_1_9_4  (
            .in0(N__3173),
            .in1(N__3145),
            .in2(N__3393),
            .in3(N__3409),
            .lcout(),
            .ltout(\Instance1.un1_r_Count_10lt11_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance1.r_Count_RNID9RS4_12_LC_1_9_5 .C_ON=1'b0;
    defparam \Instance1.r_Count_RNID9RS4_12_LC_1_9_5 .SEQ_MODE=4'b0000;
    defparam \Instance1.r_Count_RNID9RS4_12_LC_1_9_5 .LUT_INIT=16'b0001001100010001;
    LogicCell40 \Instance1.r_Count_RNID9RS4_12_LC_1_9_5  (
            .in0(N__3277),
            .in1(N__3259),
            .in2(N__2997),
            .in3(N__2994),
            .lcout(),
            .ltout(\Instance1.un1_r_Count_10lt17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance1.r_State_RNIK9757_LC_1_9_6 .C_ON=1'b0;
    defparam \Instance1.r_State_RNIK9757_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \Instance1.r_State_RNIK9757_LC_1_9_6 .LUT_INIT=16'b1001111110011001;
    LogicCell40 \Instance1.r_State_RNIK9757_LC_1_9_6  (
            .in0(N__3054),
            .in1(N__3018),
            .in2(N__2988),
            .in3(N__3093),
            .lcout(\Instance1.r_Count12_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance1.r_State_RNO_3_LC_1_9_7 .C_ON=1'b0;
    defparam \Instance1.r_State_RNO_3_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \Instance1.r_State_RNO_3_LC_1_9_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Instance1.r_State_RNO_3_LC_1_9_7  (
            .in0(N__3174),
            .in1(N__3391),
            .in2(N__3282),
            .in3(N__3260),
            .lcout(\Instance1.r_Count13_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance1.r_Count_RNIIVNV1_17_LC_1_10_0 .C_ON=1'b0;
    defparam \Instance1.r_Count_RNIIVNV1_17_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \Instance1.r_Count_RNIIVNV1_17_LC_1_10_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Instance1.r_Count_RNIIVNV1_17_LC_1_10_0  (
            .in0(N__3493),
            .in1(N__3541),
            .in2(N__3567),
            .in3(N__3517),
            .lcout(\Instance1.un1_r_Count_10lto17_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance1.r_State_RNO_4_LC_1_10_2 .C_ON=1'b0;
    defparam \Instance1.r_State_RNO_4_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \Instance1.r_State_RNO_4_LC_1_10_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Instance1.r_State_RNO_4_LC_1_10_2  (
            .in0(N__3206),
            .in1(N__3220),
            .in2(N__3192),
            .in3(N__3350),
            .lcout(\Instance1.r_Count13_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance1.r_Count_1_LC_1_10_5 .C_ON=1'b0;
    defparam \Instance1.r_Count_1_LC_1_10_5 .SEQ_MODE=4'b1000;
    defparam \Instance1.r_Count_1_LC_1_10_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \Instance1.r_Count_1_LC_1_10_5  (
            .in0(N__3221),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3473),
            .lcout(\Instance1.r_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7081),
            .ce(),
            .sr(N__3444));
    defparam r_Switch_1_LC_1_11_0.C_ON=1'b0;
    defparam r_Switch_1_LC_1_11_0.SEQ_MODE=4'b1000;
    defparam r_Switch_1_LC_1_11_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 r_Switch_1_LC_1_11_0 (
            .in0(N__3014),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r_SwitchZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7083),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance1.r_State_RNIPV6C_LC_1_11_1 .C_ON=1'b0;
    defparam \Instance1.r_State_RNIPV6C_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \Instance1.r_State_RNIPV6C_LC_1_11_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Instance1.r_State_RNIPV6C_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__3087),
            .in2(_gnd_net_),
            .in3(N__3012),
            .lcout(click13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance1.r_State_RNO_2_LC_1_11_3 .C_ON=1'b0;
    defparam \Instance1.r_State_RNO_2_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \Instance1.r_State_RNO_2_LC_1_11_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Instance1.r_State_RNO_2_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__3565),
            .in2(_gnd_net_),
            .in3(N__3494),
            .lcout(),
            .ltout(\Instance1.r_Count13_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance1.r_State_RNO_0_LC_1_11_4 .C_ON=1'b0;
    defparam \Instance1.r_State_RNO_0_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \Instance1.r_State_RNO_0_LC_1_11_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Instance1.r_State_RNO_0_LC_1_11_4  (
            .in0(N__3471),
            .in1(N__3081),
            .in2(N__3072),
            .in3(N__3150),
            .lcout(\Instance1.r_Count13_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance1.r_State_RNO_1_LC_1_11_6 .C_ON=1'b0;
    defparam \Instance1.r_State_RNO_1_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \Instance1.r_State_RNO_1_LC_1_11_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \Instance1.r_State_RNO_1_LC_1_11_6  (
            .in0(N__3069),
            .in1(N__3303),
            .in2(N__3327),
            .in3(N__3063),
            .lcout(),
            .ltout(\Instance1.r_Count13_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance1.r_State_LC_1_11_7 .C_ON=1'b0;
    defparam \Instance1.r_State_LC_1_11_7 .SEQ_MODE=4'b1000;
    defparam \Instance1.r_State_LC_1_11_7 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \Instance1.r_State_LC_1_11_7  (
            .in0(N__3053),
            .in1(N__3027),
            .in2(N__3021),
            .in3(N__3013),
            .lcout(w_Switch_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7083),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance2.r_State_RNIHFHJ2_LC_1_12_1 .C_ON=1'b0;
    defparam \Instance2.r_State_RNIHFHJ2_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \Instance2.r_State_RNIHFHJ2_LC_1_12_1 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \Instance2.r_State_RNIHFHJ2_LC_1_12_1  (
            .in0(N__4579),
            .in1(N__3987),
            .in2(_gnd_net_),
            .in3(N__4761),
            .lcout(un1_click17_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_Switch_2_RNIK7A11_LC_1_12_2.C_ON=1'b0;
    defparam r_Switch_2_RNIK7A11_LC_1_12_2.SEQ_MODE=4'b0000;
    defparam r_Switch_2_RNIK7A11_LC_1_12_2.LUT_INIT=16'b1101110111001100;
    LogicCell40 r_Switch_2_RNIK7A11_LC_1_12_2 (
            .in0(N__4917),
            .in1(N__4578),
            .in2(_gnd_net_),
            .in3(N__4833),
            .lcout(r_Switch_2_RNIK7AZ0Z11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sevsegl_RNO_0_2_LC_1_12_5.C_ON=1'b0;
    defparam sevsegl_RNO_0_2_LC_1_12_5.SEQ_MODE=4'b0000;
    defparam sevsegl_RNO_0_2_LC_1_12_5.LUT_INIT=16'b0011001110101010;
    LogicCell40 sevsegl_RNO_0_2_LC_1_12_5 (
            .in0(N__4332),
            .in1(N__4527),
            .in2(_gnd_net_),
            .in3(N__4806),
            .lcout(),
            .ltout(sevsegl_RNO_0Z0Z_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sevsegl_2_LC_1_12_6.C_ON=1'b0;
    defparam sevsegl_2_LC_1_12_6.SEQ_MODE=4'b1000;
    defparam sevsegl_2_LC_1_12_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 sevsegl_2_LC_1_12_6 (
            .in0(_gnd_net_),
            .in1(N__3123),
            .in2(N__3126),
            .in3(N__3881),
            .lcout(sevseglZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7085),
            .ce(N__3842),
            .sr(_gnd_net_));
    defparam sevsegl_RNO_1_2_LC_1_13_0.C_ON=1'b0;
    defparam sevsegl_RNO_1_2_LC_1_13_0.SEQ_MODE=4'b0000;
    defparam sevsegl_RNO_1_2_LC_1_13_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 sevsegl_RNO_1_2_LC_1_13_0 (
            .in0(N__4710),
            .in1(N__3099),
            .in2(_gnd_net_),
            .in3(N__4604),
            .lcout(sevsegl_RNO_1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sevsegr_RNO_0_0_LC_1_13_1.C_ON=1'b0;
    defparam sevsegr_RNO_0_0_LC_1_13_1.SEQ_MODE=4'b0000;
    defparam sevsegr_RNO_0_0_LC_1_13_1.LUT_INIT=16'b0101010100101110;
    LogicCell40 sevsegr_RNO_0_0_LC_1_13_1 (
            .in0(N__4386),
            .in1(N__4809),
            .in2(N__4491),
            .in3(N__3880),
            .lcout(sevsegr_7_ns_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SegInst1.r_HexEncode_i_6_LC_1_13_2 .C_ON=1'b0;
    defparam \SegInst1.r_HexEncode_i_6_LC_1_13_2 .SEQ_MODE=4'b1000;
    defparam \SegInst1.r_HexEncode_i_6_LC_1_13_2 .LUT_INIT=16'b0110000100000010;
    LogicCell40 \SegInst1.r_HexEncode_i_6_LC_1_13_2  (
            .in0(N__6060),
            .in1(N__6017),
            .in2(N__5970),
            .in3(N__5913),
            .lcout(r_HexEncode_i_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7088),
            .ce(),
            .sr(_gnd_net_));
    defparam \SegInst2.r_HexEncode_i_1_LC_1_13_3 .C_ON=1'b0;
    defparam \SegInst2.r_HexEncode_i_1_LC_1_13_3 .SEQ_MODE=4'b1000;
    defparam \SegInst2.r_HexEncode_i_1_LC_1_13_3 .LUT_INIT=16'b0010110100000100;
    LogicCell40 \SegInst2.r_HexEncode_i_1_LC_1_13_3  (
            .in0(N__3721),
            .in1(N__3676),
            .in2(N__3651),
            .in3(N__3768),
            .lcout(r_HexEncode_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7088),
            .ce(),
            .sr(_gnd_net_));
    defparam \SegInst1.r_HexEncode_i_5_LC_1_13_4 .C_ON=1'b0;
    defparam \SegInst1.r_HexEncode_i_5_LC_1_13_4 .SEQ_MODE=4'b1000;
    defparam \SegInst1.r_HexEncode_i_5_LC_1_13_4 .LUT_INIT=16'b1100001010101000;
    LogicCell40 \SegInst1.r_HexEncode_i_5_LC_1_13_4  (
            .in0(N__6059),
            .in1(N__6016),
            .in2(N__5969),
            .in3(N__5912),
            .lcout(r_HexEncode_i_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7088),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance2.SUM_2_LC_1_13_6 .C_ON=1'b0;
    defparam \Instance2.SUM_2_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \Instance2.SUM_2_LC_1_13_6 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \Instance2.SUM_2_LC_1_13_6  (
            .in0(N__4331),
            .in1(N__4454),
            .in2(_gnd_net_),
            .in3(N__4385),
            .lcout(SUM_2),
            .ltout(SUM_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sevsegr_RNO_1_2_LC_1_13_7.C_ON=1'b0;
    defparam sevsegr_RNO_1_2_LC_1_13_7.SEQ_MODE=4'b0000;
    defparam sevsegr_RNO_1_2_LC_1_13_7.LUT_INIT=16'b1111010110100000;
    LogicCell40 sevsegr_RNO_1_2_LC_1_13_7 (
            .in0(N__4605),
            .in1(_gnd_net_),
            .in2(N__3243),
            .in3(N__3906),
            .lcout(sevsegr_RNO_1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SegInst1.r_HexEncode_iZ0Z_0_LC_1_14_0 .C_ON=1'b0;
    defparam \SegInst1.r_HexEncode_iZ0Z_0_LC_1_14_0 .SEQ_MODE=4'b1000;
    defparam \SegInst1.r_HexEncode_iZ0Z_0_LC_1_14_0 .LUT_INIT=16'b0000100100100001;
    LogicCell40 \SegInst1.r_HexEncode_iZ0Z_0_LC_1_14_0  (
            .in0(N__6066),
            .in1(N__6018),
            .in2(N__5971),
            .in3(N__5914),
            .lcout(r_HexEncode_i_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7092),
            .ce(),
            .sr(_gnd_net_));
    defparam \SegInst1.r_HexEncode_i_1_LC_1_14_5 .C_ON=1'b0;
    defparam \SegInst1.r_HexEncode_i_1_LC_1_14_5 .SEQ_MODE=4'b1000;
    defparam \SegInst1.r_HexEncode_i_1_LC_1_14_5 .LUT_INIT=16'b0010100000110010;
    LogicCell40 \SegInst1.r_HexEncode_i_1_LC_1_14_5  (
            .in0(N__5915),
            .in1(N__5963),
            .in2(N__6030),
            .in3(N__6067),
            .lcout(r_HexEncode_i_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7092),
            .ce(),
            .sr(_gnd_net_));
    defparam \SegInst2.r_HexEncode_i_6_LC_1_16_3 .C_ON=1'b0;
    defparam \SegInst2.r_HexEncode_i_6_LC_1_16_3 .SEQ_MODE=4'b1000;
    defparam \SegInst2.r_HexEncode_i_6_LC_1_16_3 .LUT_INIT=16'b0110000000010100;
    LogicCell40 \SegInst2.r_HexEncode_i_6_LC_1_16_3  (
            .in0(N__3708),
            .in1(N__3741),
            .in2(N__3780),
            .in3(N__3661),
            .lcout(r_HexEncode_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7102),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance1.r_Count_2_cry_1_c_LC_2_9_0 .C_ON=1'b1;
    defparam \Instance1.r_Count_2_cry_1_c_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \Instance1.r_Count_2_cry_1_c_LC_2_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \Instance1.r_Count_2_cry_1_c_LC_2_9_0  (
            .in0(_gnd_net_),
            .in1(N__3222),
            .in2(N__3477),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_9_0_),
            .carryout(\Instance1.r_Count_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance1.r_Count_2_LC_2_9_1 .C_ON=1'b1;
    defparam \Instance1.r_Count_2_LC_2_9_1 .SEQ_MODE=4'b1000;
    defparam \Instance1.r_Count_2_LC_2_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance1.r_Count_2_LC_2_9_1  (
            .in0(_gnd_net_),
            .in1(N__3207),
            .in2(_gnd_net_),
            .in3(N__3195),
            .lcout(\Instance1.r_CountZ0Z_2 ),
            .ltout(),
            .carryin(\Instance1.r_Count_2_cry_1 ),
            .carryout(\Instance1.r_Count_2_cry_2 ),
            .clk(N__7082),
            .ce(),
            .sr(N__3445));
    defparam \Instance1.r_Count_3_LC_2_9_2 .C_ON=1'b1;
    defparam \Instance1.r_Count_3_LC_2_9_2 .SEQ_MODE=4'b1000;
    defparam \Instance1.r_Count_3_LC_2_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance1.r_Count_3_LC_2_9_2  (
            .in0(_gnd_net_),
            .in1(N__3191),
            .in2(_gnd_net_),
            .in3(N__3177),
            .lcout(\Instance1.r_CountZ0Z_3 ),
            .ltout(),
            .carryin(\Instance1.r_Count_2_cry_2 ),
            .carryout(\Instance1.r_Count_2_cry_3 ),
            .clk(N__7082),
            .ce(),
            .sr(N__3445));
    defparam \Instance1.r_Count_4_LC_2_9_3 .C_ON=1'b1;
    defparam \Instance1.r_Count_4_LC_2_9_3 .SEQ_MODE=4'b1000;
    defparam \Instance1.r_Count_4_LC_2_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance1.r_Count_4_LC_2_9_3  (
            .in0(_gnd_net_),
            .in1(N__3172),
            .in2(_gnd_net_),
            .in3(N__3153),
            .lcout(\Instance1.r_CountZ0Z_4 ),
            .ltout(),
            .carryin(\Instance1.r_Count_2_cry_3 ),
            .carryout(\Instance1.r_Count_2_cry_4 ),
            .clk(N__7082),
            .ce(),
            .sr(N__3445));
    defparam \Instance1.r_Count_5_LC_2_9_4 .C_ON=1'b1;
    defparam \Instance1.r_Count_5_LC_2_9_4 .SEQ_MODE=4'b1000;
    defparam \Instance1.r_Count_5_LC_2_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance1.r_Count_5_LC_2_9_4  (
            .in0(_gnd_net_),
            .in1(N__3146),
            .in2(_gnd_net_),
            .in3(N__3129),
            .lcout(\Instance1.r_CountZ0Z_5 ),
            .ltout(),
            .carryin(\Instance1.r_Count_2_cry_4 ),
            .carryout(\Instance1.r_Count_2_cry_5 ),
            .clk(N__7082),
            .ce(),
            .sr(N__3445));
    defparam \Instance1.r_Count_6_LC_2_9_5 .C_ON=1'b1;
    defparam \Instance1.r_Count_6_LC_2_9_5 .SEQ_MODE=4'b1000;
    defparam \Instance1.r_Count_6_LC_2_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance1.r_Count_6_LC_2_9_5  (
            .in0(_gnd_net_),
            .in1(N__3411),
            .in2(_gnd_net_),
            .in3(N__3396),
            .lcout(\Instance1.r_CountZ0Z_6 ),
            .ltout(),
            .carryin(\Instance1.r_Count_2_cry_5 ),
            .carryout(\Instance1.r_Count_2_cry_6 ),
            .clk(N__7082),
            .ce(),
            .sr(N__3445));
    defparam \Instance1.r_Count_7_LC_2_9_6 .C_ON=1'b1;
    defparam \Instance1.r_Count_7_LC_2_9_6 .SEQ_MODE=4'b1000;
    defparam \Instance1.r_Count_7_LC_2_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance1.r_Count_7_LC_2_9_6  (
            .in0(_gnd_net_),
            .in1(N__3392),
            .in2(_gnd_net_),
            .in3(N__3372),
            .lcout(\Instance1.r_CountZ0Z_7 ),
            .ltout(),
            .carryin(\Instance1.r_Count_2_cry_6 ),
            .carryout(\Instance1.r_Count_2_cry_7 ),
            .clk(N__7082),
            .ce(),
            .sr(N__3445));
    defparam \Instance1.r_Count_8_LC_2_9_7 .C_ON=1'b1;
    defparam \Instance1.r_Count_8_LC_2_9_7 .SEQ_MODE=4'b1000;
    defparam \Instance1.r_Count_8_LC_2_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance1.r_Count_8_LC_2_9_7  (
            .in0(_gnd_net_),
            .in1(N__3369),
            .in2(_gnd_net_),
            .in3(N__3354),
            .lcout(\Instance1.r_CountZ0Z_8 ),
            .ltout(),
            .carryin(\Instance1.r_Count_2_cry_7 ),
            .carryout(\Instance1.r_Count_2_cry_8 ),
            .clk(N__7082),
            .ce(),
            .sr(N__3445));
    defparam \Instance1.r_Count_9_LC_2_10_0 .C_ON=1'b1;
    defparam \Instance1.r_Count_9_LC_2_10_0 .SEQ_MODE=4'b1000;
    defparam \Instance1.r_Count_9_LC_2_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance1.r_Count_9_LC_2_10_0  (
            .in0(_gnd_net_),
            .in1(N__3349),
            .in2(_gnd_net_),
            .in3(N__3330),
            .lcout(\Instance1.r_CountZ0Z_9 ),
            .ltout(),
            .carryin(bfn_2_10_0_),
            .carryout(\Instance1.r_Count_2_cry_9 ),
            .clk(N__7084),
            .ce(),
            .sr(N__3446));
    defparam \Instance1.r_Count_10_LC_2_10_1 .C_ON=1'b1;
    defparam \Instance1.r_Count_10_LC_2_10_1 .SEQ_MODE=4'b1000;
    defparam \Instance1.r_Count_10_LC_2_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance1.r_Count_10_LC_2_10_1  (
            .in0(_gnd_net_),
            .in1(N__3323),
            .in2(_gnd_net_),
            .in3(N__3306),
            .lcout(\Instance1.r_CountZ0Z_10 ),
            .ltout(),
            .carryin(\Instance1.r_Count_2_cry_9 ),
            .carryout(\Instance1.r_Count_2_cry_10 ),
            .clk(N__7084),
            .ce(),
            .sr(N__3446));
    defparam \Instance1.r_Count_11_LC_2_10_2 .C_ON=1'b1;
    defparam \Instance1.r_Count_11_LC_2_10_2 .SEQ_MODE=4'b1000;
    defparam \Instance1.r_Count_11_LC_2_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance1.r_Count_11_LC_2_10_2  (
            .in0(_gnd_net_),
            .in1(N__3302),
            .in2(_gnd_net_),
            .in3(N__3285),
            .lcout(\Instance1.r_CountZ0Z_11 ),
            .ltout(),
            .carryin(\Instance1.r_Count_2_cry_10 ),
            .carryout(\Instance1.r_Count_2_cry_11 ),
            .clk(N__7084),
            .ce(),
            .sr(N__3446));
    defparam \Instance1.r_Count_12_LC_2_10_3 .C_ON=1'b1;
    defparam \Instance1.r_Count_12_LC_2_10_3 .SEQ_MODE=4'b1000;
    defparam \Instance1.r_Count_12_LC_2_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance1.r_Count_12_LC_2_10_3  (
            .in0(_gnd_net_),
            .in1(N__3281),
            .in2(_gnd_net_),
            .in3(N__3264),
            .lcout(\Instance1.r_CountZ0Z_12 ),
            .ltout(),
            .carryin(\Instance1.r_Count_2_cry_11 ),
            .carryout(\Instance1.r_Count_2_cry_12 ),
            .clk(N__7084),
            .ce(),
            .sr(N__3446));
    defparam \Instance1.r_Count_13_LC_2_10_4 .C_ON=1'b1;
    defparam \Instance1.r_Count_13_LC_2_10_4 .SEQ_MODE=4'b1000;
    defparam \Instance1.r_Count_13_LC_2_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance1.r_Count_13_LC_2_10_4  (
            .in0(_gnd_net_),
            .in1(N__3261),
            .in2(_gnd_net_),
            .in3(N__3246),
            .lcout(\Instance1.r_CountZ0Z_13 ),
            .ltout(),
            .carryin(\Instance1.r_Count_2_cry_12 ),
            .carryout(\Instance1.r_Count_2_cry_13 ),
            .clk(N__7084),
            .ce(),
            .sr(N__3446));
    defparam \Instance1.r_Count_14_LC_2_10_5 .C_ON=1'b1;
    defparam \Instance1.r_Count_14_LC_2_10_5 .SEQ_MODE=4'b1000;
    defparam \Instance1.r_Count_14_LC_2_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance1.r_Count_14_LC_2_10_5  (
            .in0(_gnd_net_),
            .in1(N__3566),
            .in2(_gnd_net_),
            .in3(N__3546),
            .lcout(\Instance1.r_CountZ0Z_14 ),
            .ltout(),
            .carryin(\Instance1.r_Count_2_cry_13 ),
            .carryout(\Instance1.r_Count_2_cry_14 ),
            .clk(N__7084),
            .ce(),
            .sr(N__3446));
    defparam \Instance1.r_Count_15_LC_2_10_6 .C_ON=1'b1;
    defparam \Instance1.r_Count_15_LC_2_10_6 .SEQ_MODE=4'b1000;
    defparam \Instance1.r_Count_15_LC_2_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance1.r_Count_15_LC_2_10_6  (
            .in0(_gnd_net_),
            .in1(N__3543),
            .in2(_gnd_net_),
            .in3(N__3525),
            .lcout(\Instance1.r_CountZ0Z_15 ),
            .ltout(),
            .carryin(\Instance1.r_Count_2_cry_14 ),
            .carryout(\Instance1.r_Count_2_cry_15 ),
            .clk(N__7084),
            .ce(),
            .sr(N__3446));
    defparam \Instance1.r_Count_16_LC_2_10_7 .C_ON=1'b1;
    defparam \Instance1.r_Count_16_LC_2_10_7 .SEQ_MODE=4'b1000;
    defparam \Instance1.r_Count_16_LC_2_10_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance1.r_Count_16_LC_2_10_7  (
            .in0(_gnd_net_),
            .in1(N__3521),
            .in2(_gnd_net_),
            .in3(N__3501),
            .lcout(\Instance1.r_CountZ0Z_16 ),
            .ltout(),
            .carryin(\Instance1.r_Count_2_cry_15 ),
            .carryout(\Instance1.r_Count_2_cry_16 ),
            .clk(N__7084),
            .ce(),
            .sr(N__3446));
    defparam \Instance1.r_Count_17_LC_2_11_0 .C_ON=1'b0;
    defparam \Instance1.r_Count_17_LC_2_11_0 .SEQ_MODE=4'b1000;
    defparam \Instance1.r_Count_17_LC_2_11_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Instance1.r_Count_17_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(N__3495),
            .in2(_gnd_net_),
            .in3(N__3498),
            .lcout(\Instance1.r_CountZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7086),
            .ce(),
            .sr(N__3447));
    defparam \Instance1.r_Count_0_LC_2_11_2 .C_ON=1'b0;
    defparam \Instance1.r_Count_0_LC_2_11_2 .SEQ_MODE=4'b1000;
    defparam \Instance1.r_Count_0_LC_2_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Instance1.r_Count_0_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3472),
            .lcout(\Instance1.r_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7086),
            .ce(),
            .sr(N__3447));
    defparam \alogicunit.result_1_LC_2_12_0 .C_ON=1'b0;
    defparam \alogicunit.result_1_LC_2_12_0 .SEQ_MODE=4'b1000;
    defparam \alogicunit.result_1_LC_2_12_0 .LUT_INIT=16'b1111000011110001;
    LogicCell40 \alogicunit.result_1_LC_2_12_0  (
            .in0(N__4508),
            .in1(N__4188),
            .in2(N__4106),
            .in3(N__5147),
            .lcout(right_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7089),
            .ce(N__5405),
            .sr(_gnd_net_));
    defparam \alogicunit.result_5_LC_2_12_2 .C_ON=1'b0;
    defparam \alogicunit.result_5_LC_2_12_2 .SEQ_MODE=4'b1000;
    defparam \alogicunit.result_5_LC_2_12_2 .LUT_INIT=16'b1111000111110000;
    LogicCell40 \alogicunit.result_5_LC_2_12_2  (
            .in0(N__4509),
            .in1(N__5148),
            .in2(N__4107),
            .in3(N__4053),
            .lcout(left_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7089),
            .ce(N__5405),
            .sr(_gnd_net_));
    defparam sevsegl_RNO_1_1_LC_2_12_3.C_ON=1'b0;
    defparam sevsegl_RNO_1_1_LC_2_12_3.SEQ_MODE=4'b0000;
    defparam sevsegl_RNO_1_1_LC_2_12_3.LUT_INIT=16'b0110011011110000;
    LogicCell40 sevsegl_RNO_1_1_LC_2_12_3 (
            .in0(N__4388),
            .in1(N__4460),
            .in2(N__3429),
            .in3(N__4580),
            .lcout(sevsegl_RNO_1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sevsegr_RNO_1_1_LC_2_12_4.C_ON=1'b0;
    defparam sevsegr_RNO_1_1_LC_2_12_4.SEQ_MODE=4'b0000;
    defparam sevsegr_RNO_1_1_LC_2_12_4.LUT_INIT=16'b0111001011011000;
    LogicCell40 sevsegr_RNO_1_1_LC_2_12_4 (
            .in0(N__4581),
            .in1(N__4459),
            .in2(N__3420),
            .in3(N__4387),
            .lcout(sevsegr_RNO_1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sevsegl_RNO_1_3_LC_2_12_5.C_ON=1'b0;
    defparam sevsegl_RNO_1_3_LC_2_12_5.SEQ_MODE=4'b0000;
    defparam sevsegl_RNO_1_3_LC_2_12_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 sevsegl_RNO_1_3_LC_2_12_5 (
            .in0(N__4017),
            .in1(N__3936),
            .in2(_gnd_net_),
            .in3(N__4582),
            .lcout(sevsegl_RNO_1Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sevsegr_RNO_0_3_LC_2_12_6.C_ON=1'b0;
    defparam sevsegr_RNO_0_3_LC_2_12_6.SEQ_MODE=4'b0000;
    defparam sevsegr_RNO_0_3_LC_2_12_6.LUT_INIT=16'b0111001001010000;
    LogicCell40 sevsegr_RNO_0_3_LC_2_12_6 (
            .in0(N__4807),
            .in1(N__5337),
            .in2(N__4242),
            .in3(N__5146),
            .lcout(sevsegr_RNO_0Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sevsegl_RNO_0_0_LC_2_12_7.C_ON=1'b0;
    defparam sevsegl_RNO_0_0_LC_2_12_7.SEQ_MODE=4'b0000;
    defparam sevsegl_RNO_0_0_LC_2_12_7.LUT_INIT=16'b0101010100101110;
    LogicCell40 sevsegl_RNO_0_0_LC_2_12_7 (
            .in0(N__4389),
            .in1(N__4808),
            .in2(N__4490),
            .in3(N__3879),
            .lcout(sevsegl_7_ns_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sevsegl_3_LC_2_13_0.C_ON=1'b0;
    defparam sevsegl_3_LC_2_13_0.SEQ_MODE=4'b1000;
    defparam sevsegl_3_LC_2_13_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 sevsegl_3_LC_2_13_0 (
            .in0(N__3884),
            .in1(N__4197),
            .in2(_gnd_net_),
            .in3(N__3612),
            .lcout(sevseglZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7093),
            .ce(N__3846),
            .sr(_gnd_net_));
    defparam sevsegr_1_LC_2_13_1.C_ON=1'b0;
    defparam sevsegr_1_LC_2_13_1.SEQ_MODE=4'b1000;
    defparam sevsegr_1_LC_2_13_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 sevsegr_1_LC_2_13_1 (
            .in0(N__3606),
            .in1(N__4275),
            .in2(_gnd_net_),
            .in3(N__3886),
            .lcout(sevsegrZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7093),
            .ce(N__3846),
            .sr(_gnd_net_));
    defparam sevsegr_2_LC_2_13_2.C_ON=1'b0;
    defparam sevsegr_2_LC_2_13_2.SEQ_MODE=4'b1000;
    defparam sevsegr_2_LC_2_13_2.LUT_INIT=16'b1111010110100000;
    LogicCell40 sevsegr_2_LC_2_13_2 (
            .in0(N__3887),
            .in1(_gnd_net_),
            .in2(N__3597),
            .in3(N__3996),
            .lcout(sevsegrZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7093),
            .ce(N__3846),
            .sr(_gnd_net_));
    defparam sevsegr_3_LC_2_13_3.C_ON=1'b0;
    defparam sevsegr_3_LC_2_13_3.SEQ_MODE=4'b1000;
    defparam sevsegr_3_LC_2_13_3.LUT_INIT=16'b1100110010101010;
    LogicCell40 sevsegr_3_LC_2_13_3 (
            .in0(N__3588),
            .in1(N__3918),
            .in2(_gnd_net_),
            .in3(N__3888),
            .lcout(sevsegrZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7093),
            .ce(N__3846),
            .sr(_gnd_net_));
    defparam sevsegl_1_LC_2_13_4.C_ON=1'b0;
    defparam sevsegl_1_LC_2_13_4.SEQ_MODE=4'b1000;
    defparam sevsegl_1_LC_2_13_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 sevsegl_1_LC_2_13_4 (
            .in0(N__3883),
            .in1(N__3579),
            .in2(_gnd_net_),
            .in3(N__4251),
            .lcout(sevseglZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7093),
            .ce(N__3846),
            .sr(_gnd_net_));
    defparam sevsegr_0_LC_2_13_5.C_ON=1'b0;
    defparam sevsegr_0_LC_2_13_5.SEQ_MODE=4'b1000;
    defparam sevsegr_0_LC_2_13_5.LUT_INIT=16'b1011100010101010;
    LogicCell40 sevsegr_0_LC_2_13_5 (
            .in0(N__3573),
            .in1(N__4621),
            .in2(N__3957),
            .in3(N__3885),
            .lcout(sevsegrZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7093),
            .ce(N__3846),
            .sr(_gnd_net_));
    defparam sevsegl_0_LC_2_13_7.C_ON=1'b0;
    defparam sevsegl_0_LC_2_13_7.SEQ_MODE=4'b1000;
    defparam sevsegl_0_LC_2_13_7.LUT_INIT=16'b1011100010101010;
    LogicCell40 sevsegl_0_LC_2_13_7 (
            .in0(N__3894),
            .in1(N__4620),
            .in2(N__4740),
            .in3(N__3882),
            .lcout(sevseglZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7093),
            .ce(N__3846),
            .sr(_gnd_net_));
    defparam \SegInst2.r_HexEncode_i_4_LC_2_16_2 .C_ON=1'b0;
    defparam \SegInst2.r_HexEncode_i_4_LC_2_16_2 .SEQ_MODE=4'b1000;
    defparam \SegInst2.r_HexEncode_i_4_LC_2_16_2 .LUT_INIT=16'b1100010000010000;
    LogicCell40 \SegInst2.r_HexEncode_i_4_LC_2_16_2  (
            .in0(N__3770),
            .in1(N__3739),
            .in2(N__3706),
            .in3(N__3659),
            .lcout(r_HexEncode_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7107),
            .ce(),
            .sr(_gnd_net_));
    defparam \SegInst2.r_HexEncode_i_0_LC_2_16_3 .C_ON=1'b0;
    defparam \SegInst2.r_HexEncode_i_0_LC_2_16_3 .SEQ_MODE=4'b1000;
    defparam \SegInst2.r_HexEncode_i_0_LC_2_16_3 .LUT_INIT=16'b0000100100100001;
    LogicCell40 \SegInst2.r_HexEncode_i_0_LC_2_16_3  (
            .in0(N__3736),
            .in1(N__3691),
            .in2(N__3662),
            .in3(N__3772),
            .lcout(r_HexEncode_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7107),
            .ce(),
            .sr(_gnd_net_));
    defparam \SegInst2.r_HexEncode_i_2_LC_2_16_4 .C_ON=1'b0;
    defparam \SegInst2.r_HexEncode_i_2_LC_2_16_4 .SEQ_MODE=4'b1000;
    defparam \SegInst2.r_HexEncode_i_2_LC_2_16_4 .LUT_INIT=16'b0000001010101110;
    LogicCell40 \SegInst2.r_HexEncode_i_2_LC_2_16_4  (
            .in0(N__3769),
            .in1(N__3737),
            .in2(N__3705),
            .in3(N__3655),
            .lcout(r_HexEncode_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7107),
            .ce(),
            .sr(_gnd_net_));
    defparam \SegInst2.r_HexEncode_i_3_LC_2_16_5 .C_ON=1'b0;
    defparam \SegInst2.r_HexEncode_i_3_LC_2_16_5 .SEQ_MODE=4'b1000;
    defparam \SegInst2.r_HexEncode_i_3_LC_2_16_5 .LUT_INIT=16'b1000100101000010;
    LogicCell40 \SegInst2.r_HexEncode_i_3_LC_2_16_5  (
            .in0(N__3738),
            .in1(N__3695),
            .in2(N__3663),
            .in3(N__3773),
            .lcout(r_HexEncode_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7107),
            .ce(),
            .sr(_gnd_net_));
    defparam \SegInst2.r_HexEncode_i_5_LC_2_16_6 .C_ON=1'b0;
    defparam \SegInst2.r_HexEncode_i_5_LC_2_16_6 .SEQ_MODE=4'b1000;
    defparam \SegInst2.r_HexEncode_i_5_LC_2_16_6 .LUT_INIT=16'b1110010001001000;
    LogicCell40 \SegInst2.r_HexEncode_i_5_LC_2_16_6  (
            .in0(N__3771),
            .in1(N__3740),
            .in2(N__3707),
            .in3(N__3660),
            .lcout(r_HexEncode_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7107),
            .ce(),
            .sr(_gnd_net_));
    defparam r_Count_1_LC_4_10_3.C_ON=1'b0;
    defparam r_Count_1_LC_4_10_3.SEQ_MODE=4'b1000;
    defparam r_Count_1_LC_4_10_3.LUT_INIT=16'b0001001011110000;
    LogicCell40 r_Count_1_LC_4_10_3 (
            .in0(N__4362),
            .in1(N__3982),
            .in2(N__4438),
            .in3(N__4623),
            .lcout(r_CountZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7090),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance2.SUM_3_LC_4_10_4 .C_ON=1'b0;
    defparam \Instance2.SUM_3_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \Instance2.SUM_3_LC_4_10_4 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \Instance2.SUM_3_LC_4_10_4  (
            .in0(N__4322),
            .in1(N__4419),
            .in2(N__4230),
            .in3(N__4359),
            .lcout(SUM_3),
            .ltout(SUM_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_Count_3_LC_4_10_5.C_ON=1'b0;
    defparam r_Count_3_LC_4_10_5.SEQ_MODE=4'b1000;
    defparam r_Count_3_LC_4_10_5.LUT_INIT=16'b0101000011001100;
    LogicCell40 r_Count_3_LC_4_10_5 (
            .in0(N__3983),
            .in1(N__4223),
            .in2(N__3615),
            .in3(N__4624),
            .lcout(r_CountZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7090),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance2.r_Count11_LC_4_10_6 .C_ON=1'b0;
    defparam \Instance2.r_Count11_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \Instance2.r_Count11_LC_4_10_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Instance2.r_Count11_LC_4_10_6  (
            .in0(N__4323),
            .in1(N__4418),
            .in2(N__4231),
            .in3(N__4360),
            .lcout(r_Count11),
            .ltout(r_Count11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_Count_0_LC_4_10_7.C_ON=1'b0;
    defparam r_Count_0_LC_4_10_7.SEQ_MODE=4'b1000;
    defparam r_Count_0_LC_4_10_7.LUT_INIT=16'b0000010110101010;
    LogicCell40 r_Count_0_LC_4_10_7 (
            .in0(N__4361),
            .in1(_gnd_net_),
            .in2(N__3963),
            .in3(N__4622),
            .lcout(r_CountZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7090),
            .ce(),
            .sr(_gnd_net_));
    defparam \alogicunit.result_13_iv_3_140_i_a4_1_LC_4_11_0 .C_ON=1'b0;
    defparam \alogicunit.result_13_iv_3_140_i_a4_1_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \alogicunit.result_13_iv_3_140_i_a4_1_LC_4_11_0 .LUT_INIT=16'b0101000001000101;
    LogicCell40 \alogicunit.result_13_iv_3_140_i_a4_1_LC_4_11_0  (
            .in0(N__5143),
            .in1(N__5327),
            .in2(N__5234),
            .in3(N__5038),
            .lcout(\alogicunit.N_95_1 ),
            .ltout(\alogicunit.N_95_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \alogicunit.result_0_LC_4_11_1 .C_ON=1'b0;
    defparam \alogicunit.result_0_LC_4_11_1 .SEQ_MODE=4'b1000;
    defparam \alogicunit.result_0_LC_4_11_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \alogicunit.result_0_LC_4_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3960),
            .in3(N__4643),
            .lcout(right_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7094),
            .ce(N__5406),
            .sr(_gnd_net_));
    defparam \alogicunit.result_3_LC_4_11_2 .C_ON=1'b0;
    defparam \alogicunit.result_3_LC_4_11_2 .SEQ_MODE=4'b1000;
    defparam \alogicunit.result_3_LC_4_11_2 .LUT_INIT=16'b1111010011111000;
    LogicCell40 \alogicunit.result_3_LC_4_11_2  (
            .in0(N__4133),
            .in1(N__4037),
            .in2(N__4647),
            .in3(N__4065),
            .lcout(right_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7094),
            .ce(N__5406),
            .sr(_gnd_net_));
    defparam sevsegr_RNO_1_3_LC_4_11_3.C_ON=1'b0;
    defparam sevsegr_RNO_1_3_LC_4_11_3.SEQ_MODE=4'b0000;
    defparam sevsegr_RNO_1_3_LC_4_11_3.LUT_INIT=16'b1110111001000100;
    LogicCell40 sevsegr_RNO_1_3_LC_4_11_3 (
            .in0(N__4606),
            .in1(N__3942),
            .in2(_gnd_net_),
            .in3(N__3929),
            .lcout(sevsegr_RNO_1Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \alogicunit.result_2_LC_4_11_4 .C_ON=1'b0;
    defparam \alogicunit.result_2_LC_4_11_4 .SEQ_MODE=4'b1000;
    defparam \alogicunit.result_2_LC_4_11_4 .LUT_INIT=16'b1010111011101010;
    LogicCell40 \alogicunit.result_2_LC_4_11_4  (
            .in0(N__4539),
            .in1(N__4036),
            .in2(N__4077),
            .in3(N__4183),
            .lcout(right_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7094),
            .ce(N__5406),
            .sr(_gnd_net_));
    defparam \alogicunit.negative_e_LC_4_11_6 .C_ON=1'b0;
    defparam \alogicunit.negative_e_LC_4_11_6 .SEQ_MODE=4'b1000;
    defparam \alogicunit.negative_e_LC_4_11_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \alogicunit.negative_e_LC_4_11_6  (
            .in0(N__5144),
            .in1(N__5328),
            .in2(N__5235),
            .in3(N__5039),
            .lcout(negative),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7094),
            .ce(N__5406),
            .sr(_gnd_net_));
    defparam \alogicunit.un1_a_1_cry_1_c_LC_4_12_0 .C_ON=1'b1;
    defparam \alogicunit.un1_a_1_cry_1_c_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \alogicunit.un1_a_1_cry_1_c_LC_4_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \alogicunit.un1_a_1_cry_1_c_LC_4_12_0  (
            .in0(_gnd_net_),
            .in1(N__4697),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_12_0_),
            .carryout(\alogicunit.un1_a_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \alogicunit.un1_a_1_cry_1_THRU_LUT4_0_LC_4_12_1 .C_ON=1'b1;
    defparam \alogicunit.un1_a_1_cry_1_THRU_LUT4_0_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \alogicunit.un1_a_1_cry_1_THRU_LUT4_0_LC_4_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \alogicunit.un1_a_1_cry_1_THRU_LUT4_0_LC_4_12_1  (
            .in0(_gnd_net_),
            .in1(N__4178),
            .in2(_gnd_net_),
            .in3(N__4068),
            .lcout(\alogicunit.un1_a_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\alogicunit.un1_a_1_cry_1 ),
            .carryout(\alogicunit.un1_a_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \alogicunit.un1_a_1_cry_2_THRU_LUT4_0_LC_4_12_2 .C_ON=1'b1;
    defparam \alogicunit.un1_a_1_cry_2_THRU_LUT4_0_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \alogicunit.un1_a_1_cry_2_THRU_LUT4_0_LC_4_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \alogicunit.un1_a_1_cry_2_THRU_LUT4_0_LC_4_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4134),
            .in3(N__4059),
            .lcout(\alogicunit.un1_a_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\alogicunit.un1_a_1_cry_2 ),
            .carryout(\alogicunit.un1_a_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \alogicunit.result_RNO_0_4_LC_4_12_3 .C_ON=1'b1;
    defparam \alogicunit.result_RNO_0_4_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \alogicunit.result_RNO_0_4_LC_4_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \alogicunit.result_RNO_0_4_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(N__5363),
            .in2(N__4008),
            .in3(N__4056),
            .lcout(\alogicunit.result_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\alogicunit.un1_a_1_cry_3 ),
            .carryout(\alogicunit.un1_a_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \alogicunit.result_RNO_0_5_LC_4_12_4 .C_ON=1'b1;
    defparam \alogicunit.result_RNO_0_5_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \alogicunit.result_RNO_0_5_LC_4_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \alogicunit.result_RNO_0_5_LC_4_12_4  (
            .in0(_gnd_net_),
            .in1(N__6105),
            .in2(N__4187),
            .in3(N__4044),
            .lcout(\alogicunit.result_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\alogicunit.un1_a_1_cry_4 ),
            .carryout(\alogicunit.un1_a_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \alogicunit.result_RNO_0_6_LC_4_12_5 .C_ON=1'b1;
    defparam \alogicunit.result_RNO_0_6_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \alogicunit.result_RNO_0_6_LC_4_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \alogicunit.result_RNO_0_6_LC_4_12_5  (
            .in0(_gnd_net_),
            .in1(N__5364),
            .in2(N__4260),
            .in3(N__4041),
            .lcout(\alogicunit.result_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\alogicunit.un1_a_1_cry_5 ),
            .carryout(\alogicunit.un1_a_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \alogicunit.result_7_LC_4_12_6 .C_ON=1'b0;
    defparam \alogicunit.result_7_LC_4_12_6 .SEQ_MODE=4'b1000;
    defparam \alogicunit.result_7_LC_4_12_6 .LUT_INIT=16'b1101110011101100;
    LogicCell40 \alogicunit.result_7_LC_4_12_6  (
            .in0(N__4182),
            .in1(N__4538),
            .in2(N__4038),
            .in3(N__4020),
            .lcout(left_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7098),
            .ce(N__5404),
            .sr(_gnd_net_));
    defparam \alogicunit.m26_l_fx_0_LC_4_13_0 .C_ON=1'b0;
    defparam \alogicunit.m26_l_fx_0_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \alogicunit.m26_l_fx_0_LC_4_13_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \alogicunit.m26_l_fx_0_LC_4_13_0  (
            .in0(_gnd_net_),
            .in1(N__5356),
            .in2(_gnd_net_),
            .in3(N__4160),
            .lcout(\alogicunit.m26_l_fxZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance2.un1_w_Switch_3_1_LC_4_13_1 .C_ON=1'b0;
    defparam \Instance2.un1_w_Switch_3_1_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \Instance2.un1_w_Switch_3_1_LC_4_13_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Instance2.un1_w_Switch_3_1_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(N__6555),
            .in2(_gnd_net_),
            .in3(N__4266),
            .lcout(un1_click13_1_sn),
            .ltout(un1_click13_1_sn_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sevsegr_RNO_0_2_LC_4_13_2.C_ON=1'b0;
    defparam sevsegr_RNO_0_2_LC_4_13_2.SEQ_MODE=4'b0000;
    defparam sevsegr_RNO_0_2_LC_4_13_2.LUT_INIT=16'b0000110011111100;
    LogicCell40 sevsegr_RNO_0_2_LC_4_13_2 (
            .in0(_gnd_net_),
            .in1(N__4327),
            .in2(N__3999),
            .in3(N__4520),
            .lcout(sevsegr_RNO_0Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sevsegr_RNO_0_1_LC_4_13_3.C_ON=1'b0;
    defparam sevsegr_RNO_0_1_LC_4_13_3.SEQ_MODE=4'b0000;
    defparam sevsegr_RNO_0_1_LC_4_13_3.LUT_INIT=16'b1111110010101100;
    LogicCell40 sevsegr_RNO_0_1_LC_4_13_3 (
            .in0(N__5024),
            .in1(N__4455),
            .in2(N__4805),
            .in3(N__4086),
            .lcout(sevsegr_RNO_0Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_Switch_3_LC_4_13_4.C_ON=1'b0;
    defparam r_Switch_3_LC_4_13_4.SEQ_MODE=4'b1000;
    defparam r_Switch_3_LC_4_13_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 r_Switch_3_LC_4_13_4 (
            .in0(N__6556),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r_SwitchZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7103),
            .ce(),
            .sr(_gnd_net_));
    defparam \alogicunit.m26_l_fx_LC_4_13_5 .C_ON=1'b0;
    defparam \alogicunit.m26_l_fx_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \alogicunit.m26_l_fx_LC_4_13_5 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \alogicunit.m26_l_fx_LC_4_13_5  (
            .in0(N__5357),
            .in1(_gnd_net_),
            .in2(N__4177),
            .in3(_gnd_net_),
            .lcout(\alogicunit.m26_l_fxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sevsegl_RNO_0_1_LC_4_13_6.C_ON=1'b0;
    defparam sevsegl_RNO_0_1_LC_4_13_6.SEQ_MODE=4'b0000;
    defparam sevsegl_RNO_0_1_LC_4_13_6.LUT_INIT=16'b1111110010111000;
    LogicCell40 sevsegl_RNO_0_1_LC_4_13_6 (
            .in0(N__4085),
            .in1(N__4789),
            .in2(N__4461),
            .in3(N__5025),
            .lcout(sevsegl_RNO_0Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sevsegl_RNO_0_3_LC_4_13_7.C_ON=1'b0;
    defparam sevsegl_RNO_0_3_LC_4_13_7.SEQ_MODE=4'b0000;
    defparam sevsegl_RNO_0_3_LC_4_13_7.LUT_INIT=16'b0111001001010000;
    LogicCell40 sevsegl_RNO_0_3_LC_4_13_7 (
            .in0(N__4790),
            .in1(N__5315),
            .in2(N__4238),
            .in3(N__5130),
            .lcout(sevsegl_RNO_0Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \alogicunit.m26_LC_4_14_0 .C_ON=1'b0;
    defparam \alogicunit.m26_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \alogicunit.m26_LC_4_14_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \alogicunit.m26_LC_4_14_0  (
            .in0(N__5102),
            .in1(N__5018),
            .in2(N__5225),
            .in3(N__5296),
            .lcout(\alogicunit.result24 ),
            .ltout(\alogicunit.result24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \alogicunit.un1_a_1_cry_3_c_inv_LC_4_14_1 .C_ON=1'b0;
    defparam \alogicunit.un1_a_1_cry_3_c_inv_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \alogicunit.un1_a_1_cry_3_c_inv_LC_4_14_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \alogicunit.un1_a_1_cry_3_c_inv_LC_4_14_1  (
            .in0(N__4129),
            .in1(_gnd_net_),
            .in2(N__4137),
            .in3(_gnd_net_),
            .lcout(\alogicunit.un1_a_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \alogicunit.result_13_iv_5_56_i_o4_LC_4_14_2 .C_ON=1'b0;
    defparam \alogicunit.result_13_iv_5_56_i_o4_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \alogicunit.result_13_iv_5_56_i_o4_LC_4_14_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \alogicunit.result_13_iv_5_56_i_o4_LC_4_14_2  (
            .in0(N__5209),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5022),
            .lcout(\alogicunit.N_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cu1.track_RNIVBP9_1_LC_4_14_3 .C_ON=1'b0;
    defparam \cu1.track_RNIVBP9_1_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \cu1.track_RNIVBP9_1_LC_4_14_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \cu1.track_RNIVBP9_1_LC_4_14_3  (
            .in0(N__5107),
            .in1(N__5301),
            .in2(_gnd_net_),
            .in3(N__5208),
            .lcout(cu1_track_ns_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cu1.track_RNI9MAL_1_LC_4_14_4 .C_ON=1'b0;
    defparam \cu1.track_RNI9MAL_1_LC_4_14_4 .SEQ_MODE=4'b0000;
    defparam \cu1.track_RNI9MAL_1_LC_4_14_4 .LUT_INIT=16'b1111111100111110;
    LogicCell40 \cu1.track_RNI9MAL_1_LC_4_14_4  (
            .in0(N__5207),
            .in1(N__5106),
            .in2(N__5323),
            .in3(N__5020),
            .lcout(N_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \alogicunit.m17_LC_4_14_5 .C_ON=1'b0;
    defparam \alogicunit.m17_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \alogicunit.m17_LC_4_14_5 .LUT_INIT=16'b0100000000001010;
    LogicCell40 \alogicunit.m17_LC_4_14_5  (
            .in0(N__5021),
            .in1(N__5297),
            .in2(N__5133),
            .in3(N__5210),
            .lcout(\alogicunit.N_41 ),
            .ltout(\alogicunit.N_41_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \alogicunit.result_13_iv_2_182_i_o4_LC_4_14_6 .C_ON=1'b0;
    defparam \alogicunit.result_13_iv_2_182_i_o4_LC_4_14_6 .SEQ_MODE=4'b0000;
    defparam \alogicunit.result_13_iv_2_182_i_o4_LC_4_14_6 .LUT_INIT=16'b1111110011111000;
    LogicCell40 \alogicunit.result_13_iv_2_182_i_o4_LC_4_14_6  (
            .in0(N__5303),
            .in1(N__5111),
            .in2(N__4494),
            .in3(N__5023),
            .lcout(\alogicunit.N_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cu1.track_RNI9MAL_0_1_LC_4_14_7 .C_ON=1'b0;
    defparam \cu1.track_RNI9MAL_0_1_LC_4_14_7 .SEQ_MODE=4'b0000;
    defparam \cu1.track_RNI9MAL_0_1_LC_4_14_7 .LUT_INIT=16'b1010111010111110;
    LogicCell40 \cu1.track_RNI9MAL_0_1_LC_4_14_7  (
            .in0(N__5019),
            .in1(N__5302),
            .in2(N__5132),
            .in3(N__5206),
            .lcout(track_RNI9MAL_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_Count_e_0_2_LC_4_15_0.C_ON=1'b0;
    defparam r_Count_e_0_2_LC_4_15_0.SEQ_MODE=4'b1000;
    defparam r_Count_e_0_2_LC_4_15_0.LUT_INIT=16'b0110011011001100;
    LogicCell40 r_Count_e_0_2_LC_4_15_0 (
            .in0(N__4453),
            .in1(N__4321),
            .in2(_gnd_net_),
            .in3(N__4384),
            .lcout(r_CountZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7111),
            .ce(N__4629),
            .sr(_gnd_net_));
    defparam \Instance2.r_State_RNO_3_LC_5_10_1 .C_ON=1'b0;
    defparam \Instance2.r_State_RNO_3_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \Instance2.r_State_RNO_3_LC_5_10_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Instance2.r_State_RNO_3_LC_5_10_1  (
            .in0(N__5735),
            .in1(N__5504),
            .in2(N__5715),
            .in3(N__5568),
            .lcout(),
            .ltout(\Instance2.r_Count13_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance2.r_State_RNO_0_LC_5_10_2 .C_ON=1'b0;
    defparam \Instance2.r_State_RNO_0_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \Instance2.r_State_RNO_0_LC_5_10_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Instance2.r_State_RNO_0_LC_5_10_2  (
            .in0(N__5543),
            .in1(N__6170),
            .in2(N__4281),
            .in3(N__4635),
            .lcout(\Instance2.r_Count13_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance2.r_Count_RNIIPVO_4_LC_5_10_5 .C_ON=1'b0;
    defparam \Instance2.r_Count_RNIIPVO_4_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \Instance2.r_Count_RNIIPVO_4_LC_5_10_5 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \Instance2.r_Count_RNIIPVO_4_LC_5_10_5  (
            .in0(N__5567),
            .in1(N__5542),
            .in2(N__5505),
            .in3(N__5524),
            .lcout(),
            .ltout(\Instance2.un1_r_Count_10lt11_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance2.r_Count_RNINRGT2_12_LC_5_10_6 .C_ON=1'b0;
    defparam \Instance2.r_Count_RNINRGT2_12_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \Instance2.r_Count_RNINRGT2_12_LC_5_10_6 .LUT_INIT=16'b0001001100010001;
    LogicCell40 \Instance2.r_Count_RNINRGT2_12_LC_5_10_6  (
            .in0(N__5734),
            .in1(N__5710),
            .in2(N__4278),
            .in3(N__4668),
            .lcout(\Instance2.un1_r_Count_10lt17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance2.r_State_RNO_1_LC_5_11_0 .C_ON=1'b0;
    defparam \Instance2.r_State_RNO_1_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \Instance2.r_State_RNO_1_LC_5_11_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Instance2.r_State_RNO_1_LC_5_11_0  (
            .in0(N__4653),
            .in1(N__5759),
            .in2(N__4662),
            .in3(N__5783),
            .lcout(),
            .ltout(\Instance2.r_Count13_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance2.r_State_LC_5_11_1 .C_ON=1'b0;
    defparam \Instance2.r_State_LC_5_11_1 .SEQ_MODE=4'b1000;
    defparam \Instance2.r_State_LC_5_11_1 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \Instance2.r_State_LC_5_11_1  (
            .in0(N__4871),
            .in1(N__4677),
            .in2(N__4671),
            .in3(N__4916),
            .lcout(w_Switch_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7099),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance2.r_Count_RNIGGG81_8_LC_5_11_2 .C_ON=1'b0;
    defparam \Instance2.r_Count_RNIGGG81_8_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \Instance2.r_Count_RNIGGG81_8_LC_5_11_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Instance2.r_Count_RNIGGG81_8_LC_5_11_2  (
            .in0(N__5784),
            .in1(N__5479),
            .in2(N__5760),
            .in3(N__5800),
            .lcout(\Instance2.un1_r_Count_10lto11_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance2.r_State_RNO_5_LC_5_11_4 .C_ON=1'b0;
    defparam \Instance2.r_State_RNO_5_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \Instance2.r_State_RNO_5_LC_5_11_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Instance2.r_State_RNO_5_LC_5_11_4  (
            .in0(N__5646),
            .in1(N__5525),
            .in2(N__5670),
            .in3(N__5480),
            .lcout(\Instance2.r_Count13_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance2.r_State_RNO_4_LC_5_11_5 .C_ON=1'b0;
    defparam \Instance2.r_State_RNO_4_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \Instance2.r_State_RNO_4_LC_5_11_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Instance2.r_State_RNO_4_LC_5_11_5  (
            .in0(N__5801),
            .in1(N__5589),
            .in2(N__6143),
            .in3(N__5603),
            .lcout(\Instance2.r_Count13_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \alogicunit.result_13_iv_6_14_i_o4_LC_5_11_6 .C_ON=1'b0;
    defparam \alogicunit.result_13_iv_6_14_i_o4_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \alogicunit.result_13_iv_6_14_i_o4_LC_5_11_6 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \alogicunit.result_13_iv_6_14_i_o4_LC_5_11_6  (
            .in0(N__5227),
            .in1(N__5145),
            .in2(N__5335),
            .in3(N__5040),
            .lcout(\alogicunit.N_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance2.r_State_RNO_2_LC_5_11_7 .C_ON=1'b0;
    defparam \Instance2.r_State_RNO_2_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \Instance2.r_State_RNO_2_LC_5_11_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Instance2.r_State_RNO_2_LC_5_11_7  (
            .in0(_gnd_net_),
            .in1(N__5692),
            .in2(_gnd_net_),
            .in3(N__6188),
            .lcout(\Instance2.r_Count13_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance2.r_Count_RNIMF1O1_17_LC_5_12_0 .C_ON=1'b0;
    defparam \Instance2.r_Count_RNIMF1O1_17_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \Instance2.r_Count_RNIMF1O1_17_LC_5_12_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Instance2.r_Count_RNIMF1O1_17_LC_5_12_0  (
            .in0(N__5641),
            .in1(N__6187),
            .in2(N__5694),
            .in3(N__5665),
            .lcout(\Instance2.un1_r_Count_10lto17_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam click1_LC_5_12_1.C_ON=1'b0;
    defparam click1_LC_5_12_1.SEQ_MODE=4'b1000;
    defparam click1_LC_5_12_1.LUT_INIT=16'b1111111101000100;
    LogicCell40 click1_LC_5_12_1 (
            .in0(N__4760),
            .in1(N__4963),
            .in2(_gnd_net_),
            .in3(N__4625),
            .lcout(clickZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7104),
            .ce(),
            .sr(_gnd_net_));
    defparam \alogicunit.result_13_iv_4_98_i_o4_LC_5_12_2 .C_ON=1'b0;
    defparam \alogicunit.result_13_iv_4_98_i_o4_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \alogicunit.result_13_iv_4_98_i_o4_LC_5_12_2 .LUT_INIT=16'b0001000100100110;
    LogicCell40 \alogicunit.result_13_iv_4_98_i_o4_LC_5_12_2  (
            .in0(N__5226),
            .in1(N__5142),
            .in2(N__5336),
            .in3(N__5037),
            .lcout(\alogicunit.N_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_Switch_2_LC_5_12_3.C_ON=1'b0;
    defparam r_Switch_2_LC_5_12_3.SEQ_MODE=4'b1000;
    defparam r_Switch_2_LC_5_12_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 r_Switch_2_LC_5_12_3 (
            .in0(N__4902),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r_SwitchZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7104),
            .ce(),
            .sr(_gnd_net_));
    defparam r_Switch_4_LC_5_12_4.C_ON=1'b0;
    defparam r_Switch_4_LC_5_12_4.SEQ_MODE=4'b1000;
    defparam r_Switch_4_LC_5_12_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 r_Switch_4_LC_5_12_4 (
            .in0(N__6237),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r_SwitchZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7104),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance3.r_State_LC_5_12_5 .C_ON=1'b0;
    defparam \Instance3.r_State_LC_5_12_5 .SEQ_MODE=4'b1000;
    defparam \Instance3.r_State_LC_5_12_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \Instance3.r_State_LC_5_12_5  (
            .in0(N__6795),
            .in1(N__6486),
            .in2(N__6537),
            .in3(N__6560),
            .lcout(w_Switch_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7104),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance2.r_State_RNIR73L_LC_5_12_6 .C_ON=1'b0;
    defparam \Instance2.r_State_RNIR73L_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \Instance2.r_State_RNIR73L_LC_5_12_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Instance2.r_State_RNIR73L_LC_5_12_6  (
            .in0(_gnd_net_),
            .in1(N__4901),
            .in2(_gnd_net_),
            .in3(N__4829),
            .lcout(),
            .ltout(\Instance2.click14_sn_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance2.r_State_RNINFUP1_LC_5_12_7 .C_ON=1'b0;
    defparam \Instance2.r_State_RNINFUP1_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \Instance2.r_State_RNINFUP1_LC_5_12_7 .LUT_INIT=16'b0000000000001101;
    LogicCell40 \Instance2.r_State_RNINFUP1_LC_5_12_7  (
            .in0(N__4818),
            .in1(N__6236),
            .in2(N__4812),
            .in3(N__4781),
            .lcout(Instance2_un1_click13_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \alogicunit.result_4_LC_5_13_0 .C_ON=1'b0;
    defparam \alogicunit.result_4_LC_5_13_0 .SEQ_MODE=4'b1000;
    defparam \alogicunit.result_4_LC_5_13_0 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \alogicunit.result_4_LC_5_13_0  (
            .in0(N__4685),
            .in1(N__4724),
            .in2(_gnd_net_),
            .in3(N__4746),
            .lcout(left_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7108),
            .ce(N__5400),
            .sr(_gnd_net_));
    defparam \alogicunit.result_6_LC_5_13_1 .C_ON=1'b0;
    defparam \alogicunit.result_6_LC_5_13_1 .SEQ_MODE=4'b1000;
    defparam \alogicunit.result_6_LC_5_13_1 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \alogicunit.result_6_LC_5_13_1  (
            .in0(N__4725),
            .in1(N__4686),
            .in2(_gnd_net_),
            .in3(N__4716),
            .lcout(left_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7108),
            .ce(N__5400),
            .sr(_gnd_net_));
    defparam \alogicunit.un1_a_1_cry_1_c_inv_LC_5_13_4 .C_ON=1'b0;
    defparam \alogicunit.un1_a_1_cry_1_c_inv_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \alogicunit.un1_a_1_cry_1_c_inv_LC_5_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \alogicunit.un1_a_1_cry_1_c_inv_LC_5_13_4  (
            .in0(N__6098),
            .in1(N__4698),
            .in2(_gnd_net_),
            .in3(N__5355),
            .lcout(\alogicunit.un1_a_1_cry_1_c_invZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \alogicunit.result_13_iv_2_182_i_a2_LC_5_14_0 .C_ON=1'b0;
    defparam \alogicunit.result_13_iv_2_182_i_a2_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \alogicunit.result_13_iv_2_182_i_a2_LC_5_14_0 .LUT_INIT=16'b0010001000110011;
    LogicCell40 \alogicunit.result_13_iv_2_182_i_a2_LC_5_14_0  (
            .in0(N__4990),
            .in1(N__5101),
            .in2(_gnd_net_),
            .in3(N__5201),
            .lcout(\alogicunit.N_102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cu1.track_0_LC_5_14_1 .C_ON=1'b0;
    defparam \cu1.track_0_LC_5_14_1 .SEQ_MODE=4'b1000;
    defparam \cu1.track_0_LC_5_14_1 .LUT_INIT=16'b0100010001100110;
    LogicCell40 \cu1.track_0_LC_5_14_1  (
            .in0(N__4955),
            .in1(N__5295),
            .in2(_gnd_net_),
            .in3(N__4991),
            .lcout(current_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7112),
            .ce(),
            .sr(_gnd_net_));
    defparam \cu1.track_1_LC_5_14_2 .C_ON=1'b0;
    defparam \cu1.track_1_LC_5_14_2 .SEQ_MODE=4'b1000;
    defparam \cu1.track_1_LC_5_14_2 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \cu1.track_1_LC_5_14_2  (
            .in0(N__4959),
            .in1(N__5320),
            .in2(_gnd_net_),
            .in3(N__5202),
            .lcout(current_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7112),
            .ce(),
            .sr(_gnd_net_));
    defparam \cu1.track_2_LC_5_14_3 .C_ON=1'b0;
    defparam \cu1.track_2_LC_5_14_3 .SEQ_MODE=4'b1000;
    defparam \cu1.track_2_LC_5_14_3 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \cu1.track_2_LC_5_14_3  (
            .in0(N__5321),
            .in1(N__5223),
            .in2(N__4964),
            .in3(N__5118),
            .lcout(current_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7112),
            .ce(),
            .sr(_gnd_net_));
    defparam \SegInst1.r_HexEncode_i_4_LC_5_14_5 .C_ON=1'b0;
    defparam \SegInst1.r_HexEncode_i_4_LC_5_14_5 .SEQ_MODE=4'b1000;
    defparam \SegInst1.r_HexEncode_i_4_LC_5_14_5 .LUT_INIT=16'b1000000010100100;
    LogicCell40 \SegInst1.r_HexEncode_i_4_LC_5_14_5  (
            .in0(N__6078),
            .in1(N__6031),
            .in2(N__5989),
            .in3(N__5927),
            .lcout(r_HexEncode_i_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7112),
            .ce(),
            .sr(_gnd_net_));
    defparam \alogicunit.m34_LC_5_14_6 .C_ON=1'b0;
    defparam \alogicunit.m34_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \alogicunit.m34_LC_5_14_6 .LUT_INIT=16'b0101010101010111;
    LogicCell40 \alogicunit.m34_LC_5_14_6  (
            .in0(N__4989),
            .in1(N__5319),
            .in2(N__5141),
            .in3(N__5200),
            .lcout(\alogicunit.N_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \alogicunit.result24_i_LC_5_14_7 .C_ON=1'b0;
    defparam \alogicunit.result24_i_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \alogicunit.result24_i_LC_5_14_7 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \alogicunit.result24_i_LC_5_14_7  (
            .in0(N__5100),
            .in1(N__4988),
            .in2(N__5224),
            .in3(N__5294),
            .lcout(\alogicunit.result24_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cu1.track_e_0_3_LC_5_15_1 .C_ON=1'b0;
    defparam \cu1.track_e_0_3_LC_5_15_1 .SEQ_MODE=4'b1000;
    defparam \cu1.track_e_0_3_LC_5_15_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \cu1.track_e_0_3_LC_5_15_1  (
            .in0(N__5322),
            .in1(N__5222),
            .in2(_gnd_net_),
            .in3(N__5131),
            .lcout(current_state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7115),
            .ce(N__4965),
            .sr(_gnd_net_));
    defparam \Instance2.r_State_RNI4PC15_LC_5_16_3 .C_ON=1'b0;
    defparam \Instance2.r_State_RNI4PC15_LC_5_16_3 .SEQ_MODE=4'b0000;
    defparam \Instance2.r_State_RNI4PC15_LC_5_16_3 .LUT_INIT=16'b1100001111101011;
    LogicCell40 \Instance2.r_State_RNI4PC15_LC_5_16_3  (
            .in0(N__4926),
            .in1(N__4915),
            .in2(N__4878),
            .in3(N__4848),
            .lcout(\Instance2.r_Count12_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance4.r_Count_1_LC_6_6_0 .C_ON=1'b0;
    defparam \Instance4.r_Count_1_LC_6_6_0 .SEQ_MODE=4'b1000;
    defparam \Instance4.r_Count_1_LC_6_6_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \Instance4.r_Count_1_LC_6_6_0  (
            .in0(N__6455),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5883),
            .lcout(\Instance4.r_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7101),
            .ce(),
            .sr(N__5619));
    defparam \Instance4.r_Count_0_LC_6_6_1 .C_ON=1'b0;
    defparam \Instance4.r_Count_0_LC_6_6_1 .SEQ_MODE=4'b1000;
    defparam \Instance4.r_Count_0_LC_6_6_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Instance4.r_Count_0_LC_6_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6454),
            .lcout(\Instance4.r_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7101),
            .ce(),
            .sr(N__5619));
    defparam \Instance4.r_Count_2_cry_1_c_LC_6_7_0 .C_ON=1'b1;
    defparam \Instance4.r_Count_2_cry_1_c_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \Instance4.r_Count_2_cry_1_c_LC_6_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \Instance4.r_Count_2_cry_1_c_LC_6_7_0  (
            .in0(_gnd_net_),
            .in1(N__5882),
            .in2(N__6456),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_7_0_),
            .carryout(\Instance4.r_Count_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance4.r_Count_2_LC_6_7_1 .C_ON=1'b1;
    defparam \Instance4.r_Count_2_LC_6_7_1 .SEQ_MODE=4'b1000;
    defparam \Instance4.r_Count_2_LC_6_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance4.r_Count_2_LC_6_7_1  (
            .in0(_gnd_net_),
            .in1(N__5865),
            .in2(_gnd_net_),
            .in3(N__5436),
            .lcout(\Instance4.r_CountZ0Z_2 ),
            .ltout(),
            .carryin(\Instance4.r_Count_2_cry_1 ),
            .carryout(\Instance4.r_Count_2_cry_2 ),
            .clk(N__7095),
            .ce(),
            .sr(N__5620));
    defparam \Instance4.r_Count_3_LC_6_7_2 .C_ON=1'b1;
    defparam \Instance4.r_Count_3_LC_6_7_2 .SEQ_MODE=4'b1000;
    defparam \Instance4.r_Count_3_LC_6_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance4.r_Count_3_LC_6_7_2  (
            .in0(_gnd_net_),
            .in1(N__5852),
            .in2(_gnd_net_),
            .in3(N__5433),
            .lcout(\Instance4.r_CountZ0Z_3 ),
            .ltout(),
            .carryin(\Instance4.r_Count_2_cry_2 ),
            .carryout(\Instance4.r_Count_2_cry_3 ),
            .clk(N__7095),
            .ce(),
            .sr(N__5620));
    defparam \Instance4.r_Count_4_LC_6_7_3 .C_ON=1'b1;
    defparam \Instance4.r_Count_4_LC_6_7_3 .SEQ_MODE=4'b1000;
    defparam \Instance4.r_Count_4_LC_6_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance4.r_Count_4_LC_6_7_3  (
            .in0(_gnd_net_),
            .in1(N__5838),
            .in2(_gnd_net_),
            .in3(N__5430),
            .lcout(\Instance4.r_CountZ0Z_4 ),
            .ltout(),
            .carryin(\Instance4.r_Count_2_cry_3 ),
            .carryout(\Instance4.r_Count_2_cry_4 ),
            .clk(N__7095),
            .ce(),
            .sr(N__5620));
    defparam \Instance4.r_Count_5_LC_6_7_4 .C_ON=1'b1;
    defparam \Instance4.r_Count_5_LC_6_7_4 .SEQ_MODE=4'b1000;
    defparam \Instance4.r_Count_5_LC_6_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance4.r_Count_5_LC_6_7_4  (
            .in0(_gnd_net_),
            .in1(N__6427),
            .in2(_gnd_net_),
            .in3(N__5427),
            .lcout(\Instance4.r_CountZ0Z_5 ),
            .ltout(),
            .carryin(\Instance4.r_Count_2_cry_4 ),
            .carryout(\Instance4.r_Count_2_cry_5 ),
            .clk(N__7095),
            .ce(),
            .sr(N__5620));
    defparam \Instance4.r_Count_6_LC_6_7_5 .C_ON=1'b1;
    defparam \Instance4.r_Count_6_LC_6_7_5 .SEQ_MODE=4'b1000;
    defparam \Instance4.r_Count_6_LC_6_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance4.r_Count_6_LC_6_7_5  (
            .in0(_gnd_net_),
            .in1(N__6594),
            .in2(_gnd_net_),
            .in3(N__5424),
            .lcout(\Instance4.r_CountZ0Z_6 ),
            .ltout(),
            .carryin(\Instance4.r_Count_2_cry_5 ),
            .carryout(\Instance4.r_Count_2_cry_6 ),
            .clk(N__7095),
            .ce(),
            .sr(N__5620));
    defparam \Instance4.r_Count_7_LC_6_7_6 .C_ON=1'b1;
    defparam \Instance4.r_Count_7_LC_6_7_6 .SEQ_MODE=4'b1000;
    defparam \Instance4.r_Count_7_LC_6_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance4.r_Count_7_LC_6_7_6  (
            .in0(_gnd_net_),
            .in1(N__5819),
            .in2(_gnd_net_),
            .in3(N__5421),
            .lcout(\Instance4.r_CountZ0Z_7 ),
            .ltout(),
            .carryin(\Instance4.r_Count_2_cry_6 ),
            .carryout(\Instance4.r_Count_2_cry_7 ),
            .clk(N__7095),
            .ce(),
            .sr(N__5620));
    defparam \Instance4.r_Count_8_LC_6_7_7 .C_ON=1'b1;
    defparam \Instance4.r_Count_8_LC_6_7_7 .SEQ_MODE=4'b1000;
    defparam \Instance4.r_Count_8_LC_6_7_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance4.r_Count_8_LC_6_7_7  (
            .in0(_gnd_net_),
            .in1(N__6647),
            .in2(_gnd_net_),
            .in3(N__5418),
            .lcout(\Instance4.r_CountZ0Z_8 ),
            .ltout(),
            .carryin(\Instance4.r_Count_2_cry_7 ),
            .carryout(\Instance4.r_Count_2_cry_8 ),
            .clk(N__7095),
            .ce(),
            .sr(N__5620));
    defparam \Instance4.r_Count_9_LC_6_8_0 .C_ON=1'b1;
    defparam \Instance4.r_Count_9_LC_6_8_0 .SEQ_MODE=4'b1000;
    defparam \Instance4.r_Count_9_LC_6_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance4.r_Count_9_LC_6_8_0  (
            .in0(_gnd_net_),
            .in1(N__6318),
            .in2(_gnd_net_),
            .in3(N__5463),
            .lcout(\Instance4.r_CountZ0Z_9 ),
            .ltout(),
            .carryin(bfn_6_8_0_),
            .carryout(\Instance4.r_Count_2_cry_9 ),
            .clk(N__7087),
            .ce(),
            .sr(N__5621));
    defparam \Instance4.r_Count_10_LC_6_8_1 .C_ON=1'b1;
    defparam \Instance4.r_Count_10_LC_6_8_1 .SEQ_MODE=4'b1000;
    defparam \Instance4.r_Count_10_LC_6_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance4.r_Count_10_LC_6_8_1  (
            .in0(_gnd_net_),
            .in1(N__6335),
            .in2(_gnd_net_),
            .in3(N__5460),
            .lcout(\Instance4.r_CountZ0Z_10 ),
            .ltout(),
            .carryin(\Instance4.r_Count_2_cry_9 ),
            .carryout(\Instance4.r_Count_2_cry_10 ),
            .clk(N__7087),
            .ce(),
            .sr(N__5621));
    defparam \Instance4.r_Count_11_LC_6_8_2 .C_ON=1'b1;
    defparam \Instance4.r_Count_11_LC_6_8_2 .SEQ_MODE=4'b1000;
    defparam \Instance4.r_Count_11_LC_6_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance4.r_Count_11_LC_6_8_2  (
            .in0(_gnd_net_),
            .in1(N__6351),
            .in2(_gnd_net_),
            .in3(N__5457),
            .lcout(\Instance4.r_CountZ0Z_11 ),
            .ltout(),
            .carryin(\Instance4.r_Count_2_cry_10 ),
            .carryout(\Instance4.r_Count_2_cry_11 ),
            .clk(N__7087),
            .ce(),
            .sr(N__5621));
    defparam \Instance4.r_Count_12_LC_6_8_3 .C_ON=1'b1;
    defparam \Instance4.r_Count_12_LC_6_8_3 .SEQ_MODE=4'b1000;
    defparam \Instance4.r_Count_12_LC_6_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance4.r_Count_12_LC_6_8_3  (
            .in0(_gnd_net_),
            .in1(N__6282),
            .in2(_gnd_net_),
            .in3(N__5454),
            .lcout(\Instance4.r_CountZ0Z_12 ),
            .ltout(),
            .carryin(\Instance4.r_Count_2_cry_11 ),
            .carryout(\Instance4.r_Count_2_cry_12 ),
            .clk(N__7087),
            .ce(),
            .sr(N__5621));
    defparam \Instance4.r_Count_13_LC_6_8_4 .C_ON=1'b1;
    defparam \Instance4.r_Count_13_LC_6_8_4 .SEQ_MODE=4'b1000;
    defparam \Instance4.r_Count_13_LC_6_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance4.r_Count_13_LC_6_8_4  (
            .in0(_gnd_net_),
            .in1(N__6300),
            .in2(_gnd_net_),
            .in3(N__5451),
            .lcout(\Instance4.r_CountZ0Z_13 ),
            .ltout(),
            .carryin(\Instance4.r_Count_2_cry_12 ),
            .carryout(\Instance4.r_Count_2_cry_13 ),
            .clk(N__7087),
            .ce(),
            .sr(N__5621));
    defparam \Instance4.r_Count_14_LC_6_8_5 .C_ON=1'b1;
    defparam \Instance4.r_Count_14_LC_6_8_5 .SEQ_MODE=4'b1000;
    defparam \Instance4.r_Count_14_LC_6_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance4.r_Count_14_LC_6_8_5  (
            .in0(_gnd_net_),
            .in1(N__6389),
            .in2(_gnd_net_),
            .in3(N__5448),
            .lcout(\Instance4.r_CountZ0Z_14 ),
            .ltout(),
            .carryin(\Instance4.r_Count_2_cry_13 ),
            .carryout(\Instance4.r_Count_2_cry_14 ),
            .clk(N__7087),
            .ce(),
            .sr(N__5621));
    defparam \Instance4.r_Count_15_LC_6_8_6 .C_ON=1'b1;
    defparam \Instance4.r_Count_15_LC_6_8_6 .SEQ_MODE=4'b1000;
    defparam \Instance4.r_Count_15_LC_6_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance4.r_Count_15_LC_6_8_6  (
            .in0(_gnd_net_),
            .in1(N__6630),
            .in2(_gnd_net_),
            .in3(N__5445),
            .lcout(\Instance4.r_CountZ0Z_15 ),
            .ltout(),
            .carryin(\Instance4.r_Count_2_cry_14 ),
            .carryout(\Instance4.r_Count_2_cry_15 ),
            .clk(N__7087),
            .ce(),
            .sr(N__5621));
    defparam \Instance4.r_Count_16_LC_6_8_7 .C_ON=1'b1;
    defparam \Instance4.r_Count_16_LC_6_8_7 .SEQ_MODE=4'b1000;
    defparam \Instance4.r_Count_16_LC_6_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance4.r_Count_16_LC_6_8_7  (
            .in0(_gnd_net_),
            .in1(N__6611),
            .in2(_gnd_net_),
            .in3(N__5442),
            .lcout(\Instance4.r_CountZ0Z_16 ),
            .ltout(),
            .carryin(\Instance4.r_Count_2_cry_15 ),
            .carryout(\Instance4.r_Count_2_cry_16 ),
            .clk(N__7087),
            .ce(),
            .sr(N__5621));
    defparam \Instance4.r_Count_17_LC_6_9_0 .C_ON=1'b0;
    defparam \Instance4.r_Count_17_LC_6_9_0 .SEQ_MODE=4'b1000;
    defparam \Instance4.r_Count_17_LC_6_9_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Instance4.r_Count_17_LC_6_9_0  (
            .in0(_gnd_net_),
            .in1(N__6372),
            .in2(_gnd_net_),
            .in3(N__5439),
            .lcout(\Instance4.r_CountZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7096),
            .ce(),
            .sr(N__5622));
    defparam \Instance2.r_Count_2_cry_1_c_LC_6_10_0 .C_ON=1'b1;
    defparam \Instance2.r_Count_2_cry_1_c_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \Instance2.r_Count_2_cry_1_c_LC_6_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \Instance2.r_Count_2_cry_1_c_LC_6_10_0  (
            .in0(_gnd_net_),
            .in1(N__6144),
            .in2(N__6171),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_10_0_),
            .carryout(\Instance2.r_Count_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance2.r_Count_2_LC_6_10_1 .C_ON=1'b1;
    defparam \Instance2.r_Count_2_LC_6_10_1 .SEQ_MODE=4'b1000;
    defparam \Instance2.r_Count_2_LC_6_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance2.r_Count_2_LC_6_10_1  (
            .in0(_gnd_net_),
            .in1(N__5604),
            .in2(_gnd_net_),
            .in3(N__5592),
            .lcout(\Instance2.r_Count_0_2 ),
            .ltout(),
            .carryin(\Instance2.r_Count_2_cry_1 ),
            .carryout(\Instance2.r_Count_2_cry_2 ),
            .clk(N__7100),
            .ce(),
            .sr(N__6120));
    defparam \Instance2.r_Count_3_LC_6_10_2 .C_ON=1'b1;
    defparam \Instance2.r_Count_3_LC_6_10_2 .SEQ_MODE=4'b1000;
    defparam \Instance2.r_Count_3_LC_6_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance2.r_Count_3_LC_6_10_2  (
            .in0(_gnd_net_),
            .in1(N__5582),
            .in2(_gnd_net_),
            .in3(N__5571),
            .lcout(\Instance2.r_Count_0_3 ),
            .ltout(),
            .carryin(\Instance2.r_Count_2_cry_2 ),
            .carryout(\Instance2.r_Count_2_cry_3 ),
            .clk(N__7100),
            .ce(),
            .sr(N__6120));
    defparam \Instance2.r_Count_4_LC_6_10_3 .C_ON=1'b1;
    defparam \Instance2.r_Count_4_LC_6_10_3 .SEQ_MODE=4'b1000;
    defparam \Instance2.r_Count_4_LC_6_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance2.r_Count_4_LC_6_10_3  (
            .in0(_gnd_net_),
            .in1(N__5566),
            .in2(_gnd_net_),
            .in3(N__5547),
            .lcout(\Instance2.r_CountZ0Z_4 ),
            .ltout(),
            .carryin(\Instance2.r_Count_2_cry_3 ),
            .carryout(\Instance2.r_Count_2_cry_4 ),
            .clk(N__7100),
            .ce(),
            .sr(N__6120));
    defparam \Instance2.r_Count_5_LC_6_10_4 .C_ON=1'b1;
    defparam \Instance2.r_Count_5_LC_6_10_4 .SEQ_MODE=4'b1000;
    defparam \Instance2.r_Count_5_LC_6_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance2.r_Count_5_LC_6_10_4  (
            .in0(_gnd_net_),
            .in1(N__5544),
            .in2(_gnd_net_),
            .in3(N__5529),
            .lcout(\Instance2.r_CountZ0Z_5 ),
            .ltout(),
            .carryin(\Instance2.r_Count_2_cry_4 ),
            .carryout(\Instance2.r_Count_2_cry_5 ),
            .clk(N__7100),
            .ce(),
            .sr(N__6120));
    defparam \Instance2.r_Count_6_LC_6_10_5 .C_ON=1'b1;
    defparam \Instance2.r_Count_6_LC_6_10_5 .SEQ_MODE=4'b1000;
    defparam \Instance2.r_Count_6_LC_6_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance2.r_Count_6_LC_6_10_5  (
            .in0(_gnd_net_),
            .in1(N__5526),
            .in2(_gnd_net_),
            .in3(N__5508),
            .lcout(\Instance2.r_CountZ0Z_6 ),
            .ltout(),
            .carryin(\Instance2.r_Count_2_cry_5 ),
            .carryout(\Instance2.r_Count_2_cry_6 ),
            .clk(N__7100),
            .ce(),
            .sr(N__6120));
    defparam \Instance2.r_Count_7_LC_6_10_6 .C_ON=1'b1;
    defparam \Instance2.r_Count_7_LC_6_10_6 .SEQ_MODE=4'b1000;
    defparam \Instance2.r_Count_7_LC_6_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance2.r_Count_7_LC_6_10_6  (
            .in0(_gnd_net_),
            .in1(N__5503),
            .in2(_gnd_net_),
            .in3(N__5484),
            .lcout(\Instance2.r_CountZ0Z_7 ),
            .ltout(),
            .carryin(\Instance2.r_Count_2_cry_6 ),
            .carryout(\Instance2.r_Count_2_cry_7 ),
            .clk(N__7100),
            .ce(),
            .sr(N__6120));
    defparam \Instance2.r_Count_8_LC_6_10_7 .C_ON=1'b1;
    defparam \Instance2.r_Count_8_LC_6_10_7 .SEQ_MODE=4'b1000;
    defparam \Instance2.r_Count_8_LC_6_10_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance2.r_Count_8_LC_6_10_7  (
            .in0(_gnd_net_),
            .in1(N__5481),
            .in2(_gnd_net_),
            .in3(N__5466),
            .lcout(\Instance2.r_CountZ0Z_8 ),
            .ltout(),
            .carryin(\Instance2.r_Count_2_cry_7 ),
            .carryout(\Instance2.r_Count_2_cry_8 ),
            .clk(N__7100),
            .ce(),
            .sr(N__6120));
    defparam \Instance2.r_Count_9_LC_6_11_0 .C_ON=1'b1;
    defparam \Instance2.r_Count_9_LC_6_11_0 .SEQ_MODE=4'b1000;
    defparam \Instance2.r_Count_9_LC_6_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance2.r_Count_9_LC_6_11_0  (
            .in0(_gnd_net_),
            .in1(N__5802),
            .in2(_gnd_net_),
            .in3(N__5787),
            .lcout(\Instance2.r_CountZ0Z_9 ),
            .ltout(),
            .carryin(bfn_6_11_0_),
            .carryout(\Instance2.r_Count_2_cry_9 ),
            .clk(N__7105),
            .ce(),
            .sr(N__6119));
    defparam \Instance2.r_Count_10_LC_6_11_1 .C_ON=1'b1;
    defparam \Instance2.r_Count_10_LC_6_11_1 .SEQ_MODE=4'b1000;
    defparam \Instance2.r_Count_10_LC_6_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance2.r_Count_10_LC_6_11_1  (
            .in0(_gnd_net_),
            .in1(N__5782),
            .in2(_gnd_net_),
            .in3(N__5763),
            .lcout(\Instance2.r_CountZ0Z_10 ),
            .ltout(),
            .carryin(\Instance2.r_Count_2_cry_9 ),
            .carryout(\Instance2.r_Count_2_cry_10 ),
            .clk(N__7105),
            .ce(),
            .sr(N__6119));
    defparam \Instance2.r_Count_11_LC_6_11_2 .C_ON=1'b1;
    defparam \Instance2.r_Count_11_LC_6_11_2 .SEQ_MODE=4'b1000;
    defparam \Instance2.r_Count_11_LC_6_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance2.r_Count_11_LC_6_11_2  (
            .in0(_gnd_net_),
            .in1(N__5758),
            .in2(_gnd_net_),
            .in3(N__5739),
            .lcout(\Instance2.r_CountZ0Z_11 ),
            .ltout(),
            .carryin(\Instance2.r_Count_2_cry_10 ),
            .carryout(\Instance2.r_Count_2_cry_11 ),
            .clk(N__7105),
            .ce(),
            .sr(N__6119));
    defparam \Instance2.r_Count_12_LC_6_11_3 .C_ON=1'b1;
    defparam \Instance2.r_Count_12_LC_6_11_3 .SEQ_MODE=4'b1000;
    defparam \Instance2.r_Count_12_LC_6_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance2.r_Count_12_LC_6_11_3  (
            .in0(_gnd_net_),
            .in1(N__5736),
            .in2(_gnd_net_),
            .in3(N__5718),
            .lcout(\Instance2.r_CountZ0Z_12 ),
            .ltout(),
            .carryin(\Instance2.r_Count_2_cry_11 ),
            .carryout(\Instance2.r_Count_2_cry_12 ),
            .clk(N__7105),
            .ce(),
            .sr(N__6119));
    defparam \Instance2.r_Count_13_LC_6_11_4 .C_ON=1'b1;
    defparam \Instance2.r_Count_13_LC_6_11_4 .SEQ_MODE=4'b1000;
    defparam \Instance2.r_Count_13_LC_6_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance2.r_Count_13_LC_6_11_4  (
            .in0(_gnd_net_),
            .in1(N__5714),
            .in2(_gnd_net_),
            .in3(N__5697),
            .lcout(\Instance2.r_CountZ0Z_13 ),
            .ltout(),
            .carryin(\Instance2.r_Count_2_cry_12 ),
            .carryout(\Instance2.r_Count_2_cry_13 ),
            .clk(N__7105),
            .ce(),
            .sr(N__6119));
    defparam \Instance2.r_Count_14_LC_6_11_5 .C_ON=1'b1;
    defparam \Instance2.r_Count_14_LC_6_11_5 .SEQ_MODE=4'b1000;
    defparam \Instance2.r_Count_14_LC_6_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance2.r_Count_14_LC_6_11_5  (
            .in0(_gnd_net_),
            .in1(N__5693),
            .in2(_gnd_net_),
            .in3(N__5673),
            .lcout(\Instance2.r_CountZ0Z_14 ),
            .ltout(),
            .carryin(\Instance2.r_Count_2_cry_13 ),
            .carryout(\Instance2.r_Count_2_cry_14 ),
            .clk(N__7105),
            .ce(),
            .sr(N__6119));
    defparam \Instance2.r_Count_15_LC_6_11_6 .C_ON=1'b1;
    defparam \Instance2.r_Count_15_LC_6_11_6 .SEQ_MODE=4'b1000;
    defparam \Instance2.r_Count_15_LC_6_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance2.r_Count_15_LC_6_11_6  (
            .in0(_gnd_net_),
            .in1(N__5669),
            .in2(_gnd_net_),
            .in3(N__5649),
            .lcout(\Instance2.r_CountZ0Z_15 ),
            .ltout(),
            .carryin(\Instance2.r_Count_2_cry_14 ),
            .carryout(\Instance2.r_Count_2_cry_15 ),
            .clk(N__7105),
            .ce(),
            .sr(N__6119));
    defparam \Instance2.r_Count_16_LC_6_11_7 .C_ON=1'b1;
    defparam \Instance2.r_Count_16_LC_6_11_7 .SEQ_MODE=4'b1000;
    defparam \Instance2.r_Count_16_LC_6_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance2.r_Count_16_LC_6_11_7  (
            .in0(_gnd_net_),
            .in1(N__5645),
            .in2(_gnd_net_),
            .in3(N__5625),
            .lcout(\Instance2.r_CountZ0Z_16 ),
            .ltout(),
            .carryin(\Instance2.r_Count_2_cry_15 ),
            .carryout(\Instance2.r_Count_2_cry_16 ),
            .clk(N__7105),
            .ce(),
            .sr(N__6119));
    defparam \Instance2.r_Count_17_LC_6_12_0 .C_ON=1'b0;
    defparam \Instance2.r_Count_17_LC_6_12_0 .SEQ_MODE=4'b1000;
    defparam \Instance2.r_Count_17_LC_6_12_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Instance2.r_Count_17_LC_6_12_0  (
            .in0(_gnd_net_),
            .in1(N__6189),
            .in2(_gnd_net_),
            .in3(N__6192),
            .lcout(\Instance2.r_CountZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7109),
            .ce(),
            .sr(N__6118));
    defparam \Instance2.r_Count_0_LC_6_12_5 .C_ON=1'b0;
    defparam \Instance2.r_Count_0_LC_6_12_5 .SEQ_MODE=4'b1000;
    defparam \Instance2.r_Count_0_LC_6_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Instance2.r_Count_0_LC_6_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6165),
            .lcout(\Instance2.r_Count_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7109),
            .ce(),
            .sr(N__6118));
    defparam \Instance2.r_Count_1_LC_6_12_6 .C_ON=1'b0;
    defparam \Instance2.r_Count_1_LC_6_12_6 .SEQ_MODE=4'b1000;
    defparam \Instance2.r_Count_1_LC_6_12_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \Instance2.r_Count_1_LC_6_12_6  (
            .in0(N__6166),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6142),
            .lcout(\Instance2.r_Count_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7109),
            .ce(),
            .sr(N__6118));
    defparam CONSTANT_ONE_LUT4_LC_6_13_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_6_13_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_6_13_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_6_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SegInst1.r_HexEncode_i_3_LC_6_14_0 .C_ON=1'b0;
    defparam \SegInst1.r_HexEncode_i_3_LC_6_14_0 .SEQ_MODE=4'b1000;
    defparam \SegInst1.r_HexEncode_i_3_LC_6_14_0 .LUT_INIT=16'b1000100101000010;
    LogicCell40 \SegInst1.r_HexEncode_i_3_LC_6_14_0  (
            .in0(N__6077),
            .in1(N__6033),
            .in2(N__5991),
            .in3(N__5934),
            .lcout(r_HexEncode_i_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7116),
            .ce(),
            .sr(_gnd_net_));
    defparam \SegInst1.r_HexEncode_i_2_LC_6_14_4 .C_ON=1'b0;
    defparam \SegInst1.r_HexEncode_i_2_LC_6_14_4 .SEQ_MODE=4'b1000;
    defparam \SegInst1.r_HexEncode_i_2_LC_6_14_4 .LUT_INIT=16'b0001111100000010;
    LogicCell40 \SegInst1.r_HexEncode_i_2_LC_6_14_4  (
            .in0(N__6076),
            .in1(N__6032),
            .in2(N__5990),
            .in3(N__5933),
            .lcout(r_HexEncode_i_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7116),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance4.r_State_RNO_4_LC_7_7_1 .C_ON=1'b0;
    defparam \Instance4.r_State_RNO_4_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \Instance4.r_State_RNO_4_LC_7_7_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Instance4.r_State_RNO_4_LC_7_7_1  (
            .in0(N__5881),
            .in1(N__5864),
            .in2(N__5853),
            .in3(N__6317),
            .lcout(\Instance4.r_Count13_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance4.r_Count_RNIQHQE_4_LC_7_7_4 .C_ON=1'b0;
    defparam \Instance4.r_Count_RNIQHQE_4_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \Instance4.r_Count_RNIQHQE_4_LC_7_7_4 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \Instance4.r_Count_RNIQHQE_4_LC_7_7_4  (
            .in0(N__5818),
            .in1(N__5836),
            .in2(N__6429),
            .in3(N__6592),
            .lcout(\Instance4.un1_r_Count_10lt11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance4.r_State_RNO_3_LC_7_7_5 .C_ON=1'b0;
    defparam \Instance4.r_State_RNO_3_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \Instance4.r_State_RNO_3_LC_7_7_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Instance4.r_State_RNO_3_LC_7_7_5  (
            .in0(N__5837),
            .in1(N__6299),
            .in2(N__5823),
            .in3(N__6281),
            .lcout(),
            .ltout(\Instance4.r_Count13_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance4.r_State_RNO_0_LC_7_7_6 .C_ON=1'b0;
    defparam \Instance4.r_State_RNO_0_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \Instance4.r_State_RNO_0_LC_7_7_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Instance4.r_State_RNO_0_LC_7_7_6  (
            .in0(N__6357),
            .in1(N__6453),
            .in2(N__6432),
            .in3(N__6428),
            .lcout(\Instance4.r_Count13_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance4.r_State_RNO_1_LC_7_8_0 .C_ON=1'b0;
    defparam \Instance4.r_State_RNO_1_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \Instance4.r_State_RNO_1_LC_7_8_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Instance4.r_State_RNO_1_LC_7_8_0  (
            .in0(N__6334),
            .in1(N__6408),
            .in2(N__6576),
            .in3(N__6350),
            .lcout(),
            .ltout(\Instance4.r_Count13_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance4.r_State_LC_7_8_1 .C_ON=1'b0;
    defparam \Instance4.r_State_LC_7_8_1 .SEQ_MODE=4'b1000;
    defparam \Instance4.r_State_LC_7_8_1 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \Instance4.r_State_LC_7_8_1  (
            .in0(N__6227),
            .in1(N__6254),
            .in2(N__6402),
            .in3(N__6399),
            .lcout(w_Switch_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7091),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance4.r_Count_RNIUFK81_17_LC_7_8_2 .C_ON=1'b0;
    defparam \Instance4.r_Count_RNIUFK81_17_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \Instance4.r_Count_RNIUFK81_17_LC_7_8_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Instance4.r_Count_RNIUFK81_17_LC_7_8_2  (
            .in0(N__6370),
            .in1(N__6628),
            .in2(N__6390),
            .in3(N__6607),
            .lcout(\Instance4.un1_r_Count_10lto17_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance4.r_State_RNO_2_LC_7_8_3 .C_ON=1'b0;
    defparam \Instance4.r_State_RNO_2_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \Instance4.r_State_RNO_2_LC_7_8_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Instance4.r_State_RNO_2_LC_7_8_3  (
            .in0(_gnd_net_),
            .in1(N__6388),
            .in2(_gnd_net_),
            .in3(N__6371),
            .lcout(\Instance4.r_Count13_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance4.r_Count_RNIOCNR_8_LC_7_8_4 .C_ON=1'b0;
    defparam \Instance4.r_Count_RNIOCNR_8_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \Instance4.r_Count_RNIOCNR_8_LC_7_8_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Instance4.r_Count_RNIOCNR_8_LC_7_8_4  (
            .in0(N__6646),
            .in1(N__6349),
            .in2(N__6336),
            .in3(N__6316),
            .lcout(),
            .ltout(\Instance4.un1_r_Count_10lto11_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance4.r_Count_RNIB0SU1_12_LC_7_8_5 .C_ON=1'b0;
    defparam \Instance4.r_Count_RNIB0SU1_12_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \Instance4.r_Count_RNIB0SU1_12_LC_7_8_5 .LUT_INIT=16'b0001000101010001;
    LogicCell40 \Instance4.r_Count_RNIB0SU1_12_LC_7_8_5  (
            .in0(N__6298),
            .in1(N__6280),
            .in2(N__6264),
            .in3(N__6261),
            .lcout(),
            .ltout(\Instance4.un1_r_Count_10lt17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance4.r_State_RNI4ONP3_LC_7_8_6 .C_ON=1'b0;
    defparam \Instance4.r_State_RNI4ONP3_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \Instance4.r_State_RNI4ONP3_LC_7_8_6 .LUT_INIT=16'b1001111110011001;
    LogicCell40 \Instance4.r_State_RNI4ONP3_LC_7_8_6  (
            .in0(N__6255),
            .in1(N__6226),
            .in2(N__6213),
            .in3(N__6210),
            .lcout(\Instance4.r_Count12_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance4.r_State_RNO_5_LC_7_8_7 .C_ON=1'b0;
    defparam \Instance4.r_State_RNO_5_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \Instance4.r_State_RNO_5_LC_7_8_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Instance4.r_State_RNO_5_LC_7_8_7  (
            .in0(N__6648),
            .in1(N__6629),
            .in2(N__6612),
            .in3(N__6593),
            .lcout(\Instance4.r_Count13_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance3.r_Count_RNI1E6U3_12_LC_7_9_0 .C_ON=1'b0;
    defparam \Instance3.r_Count_RNI1E6U3_12_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \Instance3.r_Count_RNI1E6U3_12_LC_7_9_0 .LUT_INIT=16'b0001001100000011;
    LogicCell40 \Instance3.r_Count_RNI1E6U3_12_LC_7_9_0  (
            .in0(N__6474),
            .in1(N__6814),
            .in2(N__6846),
            .in3(N__6468),
            .lcout(),
            .ltout(\Instance3.un1_r_Count_10lt17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance3.r_State_RNIK8IT5_LC_7_9_1 .C_ON=1'b0;
    defparam \Instance3.r_State_RNIK8IT5_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \Instance3.r_State_RNIK8IT5_LC_7_9_1 .LUT_INIT=16'b1001111110011001;
    LogicCell40 \Instance3.r_State_RNIK8IT5_LC_7_9_1  (
            .in0(N__6567),
            .in1(N__6530),
            .in2(N__6501),
            .in3(N__6777),
            .lcout(\Instance3.r_Count12_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance3.r_State_RNO_3_LC_7_9_3 .C_ON=1'b0;
    defparam \Instance3.r_State_RNO_3_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \Instance3.r_State_RNO_3_LC_7_9_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Instance3.r_State_RNO_3_LC_7_9_3  (
            .in0(N__6841),
            .in1(N__6956),
            .in2(N__6819),
            .in3(N__6686),
            .lcout(),
            .ltout(\Instance3.r_Count13_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance3.r_State_RNO_0_LC_7_9_4 .C_ON=1'b0;
    defparam \Instance3.r_State_RNO_0_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \Instance3.r_State_RNO_0_LC_7_9_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Instance3.r_State_RNO_0_LC_7_9_4  (
            .in0(N__6668),
            .in1(N__7167),
            .in2(N__6489),
            .in3(N__6462),
            .lcout(\Instance3.r_Count13_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance3.r_Count_RNIM5TJ1_4_LC_7_9_5 .C_ON=1'b0;
    defparam \Instance3.r_Count_RNIM5TJ1_4_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \Instance3.r_Count_RNIM5TJ1_4_LC_7_9_5 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \Instance3.r_Count_RNIM5TJ1_4_LC_7_9_5  (
            .in0(N__6669),
            .in1(N__6685),
            .in2(N__6981),
            .in3(N__6955),
            .lcout(\Instance3.un1_r_Count_10lt11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance3.r_Count_RNIKU3I1_10_LC_7_9_7 .C_ON=1'b0;
    defparam \Instance3.r_Count_RNIKU3I1_10_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \Instance3.r_Count_RNIKU3I1_10_LC_7_9_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Instance3.r_Count_RNIKU3I1_10_LC_7_9_7  (
            .in0(N__6870),
            .in1(N__6937),
            .in2(N__6897),
            .in3(N__6916),
            .lcout(\Instance3.un1_r_Count_10lto11_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance3.r_State_RNO_2_LC_7_10_0 .C_ON=1'b0;
    defparam \Instance3.r_State_RNO_2_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \Instance3.r_State_RNO_2_LC_7_10_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Instance3.r_State_RNO_2_LC_7_10_0  (
            .in0(_gnd_net_),
            .in1(N__7249),
            .in2(_gnd_net_),
            .in3(N__7181),
            .lcout(\Instance3.r_Count13_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance3.r_State_RNO_4_LC_7_10_1 .C_ON=1'b0;
    defparam \Instance3.r_State_RNO_4_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \Instance3.r_State_RNO_4_LC_7_10_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Instance3.r_State_RNO_4_LC_7_10_1  (
            .in0(N__6719),
            .in1(N__7137),
            .in2(N__6705),
            .in3(N__6917),
            .lcout(),
            .ltout(\Instance3.r_Count13_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance3.r_State_RNO_1_LC_7_10_2 .C_ON=1'b0;
    defparam \Instance3.r_State_RNO_1_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \Instance3.r_State_RNO_1_LC_7_10_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Instance3.r_State_RNO_1_LC_7_10_2  (
            .in0(N__6783),
            .in1(N__6868),
            .in2(N__6798),
            .in3(N__6892),
            .lcout(\Instance3.r_Count13_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance3.r_State_RNO_5_LC_7_10_3 .C_ON=1'b0;
    defparam \Instance3.r_State_RNO_5_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \Instance3.r_State_RNO_5_LC_7_10_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Instance3.r_State_RNO_5_LC_7_10_3  (
            .in0(N__7205),
            .in1(N__6979),
            .in2(N__7230),
            .in3(N__6938),
            .lcout(\Instance3.r_Count13_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance3.r_Count_RNIQVAG1_17_LC_7_10_7 .C_ON=1'b0;
    defparam \Instance3.r_Count_RNIQVAG1_17_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \Instance3.r_Count_RNIQVAG1_17_LC_7_10_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Instance3.r_Count_RNIQVAG1_17_LC_7_10_7  (
            .in0(N__7180),
            .in1(N__7225),
            .in2(N__7251),
            .in3(N__7204),
            .lcout(\Instance3.un1_r_Count_10lto17_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_1_1_LC_8_8_4.C_ON=1'b0;
    defparam o_LED_1_1_LC_8_8_4.SEQ_MODE=4'b1000;
    defparam o_LED_1_1_LC_8_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 o_LED_1_1_LC_8_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6771),
            .lcout(o_LED_1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7097),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance3.r_Count_2_cry_1_c_LC_8_9_0 .C_ON=1'b1;
    defparam \Instance3.r_Count_2_cry_1_c_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \Instance3.r_Count_2_cry_1_c_LC_8_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \Instance3.r_Count_2_cry_1_c_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(N__7135),
            .in2(N__7163),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(\Instance3.r_Count_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Instance3.r_Count_2_LC_8_9_1 .C_ON=1'b1;
    defparam \Instance3.r_Count_2_LC_8_9_1 .SEQ_MODE=4'b1000;
    defparam \Instance3.r_Count_2_LC_8_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance3.r_Count_2_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(N__6720),
            .in2(_gnd_net_),
            .in3(N__6708),
            .lcout(\Instance3.r_CountZ0Z_2 ),
            .ltout(),
            .carryin(\Instance3.r_Count_2_cry_1 ),
            .carryout(\Instance3.r_Count_2_cry_2 ),
            .clk(N__7106),
            .ce(),
            .sr(N__6999));
    defparam \Instance3.r_Count_3_LC_8_9_2 .C_ON=1'b1;
    defparam \Instance3.r_Count_3_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \Instance3.r_Count_3_LC_8_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance3.r_Count_3_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(N__6704),
            .in2(_gnd_net_),
            .in3(N__6690),
            .lcout(\Instance3.r_CountZ0Z_3 ),
            .ltout(),
            .carryin(\Instance3.r_Count_2_cry_2 ),
            .carryout(\Instance3.r_Count_2_cry_3 ),
            .clk(N__7106),
            .ce(),
            .sr(N__6999));
    defparam \Instance3.r_Count_4_LC_8_9_3 .C_ON=1'b1;
    defparam \Instance3.r_Count_4_LC_8_9_3 .SEQ_MODE=4'b1000;
    defparam \Instance3.r_Count_4_LC_8_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance3.r_Count_4_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__6687),
            .in2(_gnd_net_),
            .in3(N__6672),
            .lcout(\Instance3.r_CountZ0Z_4 ),
            .ltout(),
            .carryin(\Instance3.r_Count_2_cry_3 ),
            .carryout(\Instance3.r_Count_2_cry_4 ),
            .clk(N__7106),
            .ce(),
            .sr(N__6999));
    defparam \Instance3.r_Count_5_LC_8_9_4 .C_ON=1'b1;
    defparam \Instance3.r_Count_5_LC_8_9_4 .SEQ_MODE=4'b1000;
    defparam \Instance3.r_Count_5_LC_8_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance3.r_Count_5_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(N__6667),
            .in2(_gnd_net_),
            .in3(N__6984),
            .lcout(\Instance3.r_CountZ0Z_5 ),
            .ltout(),
            .carryin(\Instance3.r_Count_2_cry_4 ),
            .carryout(\Instance3.r_Count_2_cry_5 ),
            .clk(N__7106),
            .ce(),
            .sr(N__6999));
    defparam \Instance3.r_Count_6_LC_8_9_5 .C_ON=1'b1;
    defparam \Instance3.r_Count_6_LC_8_9_5 .SEQ_MODE=4'b1000;
    defparam \Instance3.r_Count_6_LC_8_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance3.r_Count_6_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(N__6980),
            .in2(_gnd_net_),
            .in3(N__6960),
            .lcout(\Instance3.r_CountZ0Z_6 ),
            .ltout(),
            .carryin(\Instance3.r_Count_2_cry_5 ),
            .carryout(\Instance3.r_Count_2_cry_6 ),
            .clk(N__7106),
            .ce(),
            .sr(N__6999));
    defparam \Instance3.r_Count_7_LC_8_9_6 .C_ON=1'b1;
    defparam \Instance3.r_Count_7_LC_8_9_6 .SEQ_MODE=4'b1000;
    defparam \Instance3.r_Count_7_LC_8_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance3.r_Count_7_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(N__6957),
            .in2(_gnd_net_),
            .in3(N__6942),
            .lcout(\Instance3.r_CountZ0Z_7 ),
            .ltout(),
            .carryin(\Instance3.r_Count_2_cry_6 ),
            .carryout(\Instance3.r_Count_2_cry_7 ),
            .clk(N__7106),
            .ce(),
            .sr(N__6999));
    defparam \Instance3.r_Count_8_LC_8_9_7 .C_ON=1'b1;
    defparam \Instance3.r_Count_8_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \Instance3.r_Count_8_LC_8_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance3.r_Count_8_LC_8_9_7  (
            .in0(_gnd_net_),
            .in1(N__6939),
            .in2(_gnd_net_),
            .in3(N__6921),
            .lcout(\Instance3.r_CountZ0Z_8 ),
            .ltout(),
            .carryin(\Instance3.r_Count_2_cry_7 ),
            .carryout(\Instance3.r_Count_2_cry_8 ),
            .clk(N__7106),
            .ce(),
            .sr(N__6999));
    defparam \Instance3.r_Count_9_LC_8_10_0 .C_ON=1'b1;
    defparam \Instance3.r_Count_9_LC_8_10_0 .SEQ_MODE=4'b1000;
    defparam \Instance3.r_Count_9_LC_8_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance3.r_Count_9_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(N__6918),
            .in2(_gnd_net_),
            .in3(N__6900),
            .lcout(\Instance3.r_CountZ0Z_9 ),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(\Instance3.r_Count_2_cry_9 ),
            .clk(N__7110),
            .ce(),
            .sr(N__7001));
    defparam \Instance3.r_Count_10_LC_8_10_1 .C_ON=1'b1;
    defparam \Instance3.r_Count_10_LC_8_10_1 .SEQ_MODE=4'b1000;
    defparam \Instance3.r_Count_10_LC_8_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance3.r_Count_10_LC_8_10_1  (
            .in0(_gnd_net_),
            .in1(N__6893),
            .in2(_gnd_net_),
            .in3(N__6873),
            .lcout(\Instance3.r_CountZ0Z_10 ),
            .ltout(),
            .carryin(\Instance3.r_Count_2_cry_9 ),
            .carryout(\Instance3.r_Count_2_cry_10 ),
            .clk(N__7110),
            .ce(),
            .sr(N__7001));
    defparam \Instance3.r_Count_11_LC_8_10_2 .C_ON=1'b1;
    defparam \Instance3.r_Count_11_LC_8_10_2 .SEQ_MODE=4'b1000;
    defparam \Instance3.r_Count_11_LC_8_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance3.r_Count_11_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(N__6869),
            .in2(_gnd_net_),
            .in3(N__6849),
            .lcout(\Instance3.r_CountZ0Z_11 ),
            .ltout(),
            .carryin(\Instance3.r_Count_2_cry_10 ),
            .carryout(\Instance3.r_Count_2_cry_11 ),
            .clk(N__7110),
            .ce(),
            .sr(N__7001));
    defparam \Instance3.r_Count_12_LC_8_10_3 .C_ON=1'b1;
    defparam \Instance3.r_Count_12_LC_8_10_3 .SEQ_MODE=4'b1000;
    defparam \Instance3.r_Count_12_LC_8_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance3.r_Count_12_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(N__6842),
            .in2(_gnd_net_),
            .in3(N__6822),
            .lcout(\Instance3.r_CountZ0Z_12 ),
            .ltout(),
            .carryin(\Instance3.r_Count_2_cry_11 ),
            .carryout(\Instance3.r_Count_2_cry_12 ),
            .clk(N__7110),
            .ce(),
            .sr(N__7001));
    defparam \Instance3.r_Count_13_LC_8_10_4 .C_ON=1'b1;
    defparam \Instance3.r_Count_13_LC_8_10_4 .SEQ_MODE=4'b1000;
    defparam \Instance3.r_Count_13_LC_8_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance3.r_Count_13_LC_8_10_4  (
            .in0(_gnd_net_),
            .in1(N__6818),
            .in2(_gnd_net_),
            .in3(N__6801),
            .lcout(\Instance3.r_CountZ0Z_13 ),
            .ltout(),
            .carryin(\Instance3.r_Count_2_cry_12 ),
            .carryout(\Instance3.r_Count_2_cry_13 ),
            .clk(N__7110),
            .ce(),
            .sr(N__7001));
    defparam \Instance3.r_Count_14_LC_8_10_5 .C_ON=1'b1;
    defparam \Instance3.r_Count_14_LC_8_10_5 .SEQ_MODE=4'b1000;
    defparam \Instance3.r_Count_14_LC_8_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance3.r_Count_14_LC_8_10_5  (
            .in0(_gnd_net_),
            .in1(N__7250),
            .in2(_gnd_net_),
            .in3(N__7233),
            .lcout(\Instance3.r_CountZ0Z_14 ),
            .ltout(),
            .carryin(\Instance3.r_Count_2_cry_13 ),
            .carryout(\Instance3.r_Count_2_cry_14 ),
            .clk(N__7110),
            .ce(),
            .sr(N__7001));
    defparam \Instance3.r_Count_15_LC_8_10_6 .C_ON=1'b1;
    defparam \Instance3.r_Count_15_LC_8_10_6 .SEQ_MODE=4'b1000;
    defparam \Instance3.r_Count_15_LC_8_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance3.r_Count_15_LC_8_10_6  (
            .in0(_gnd_net_),
            .in1(N__7229),
            .in2(_gnd_net_),
            .in3(N__7209),
            .lcout(\Instance3.r_CountZ0Z_15 ),
            .ltout(),
            .carryin(\Instance3.r_Count_2_cry_14 ),
            .carryout(\Instance3.r_Count_2_cry_15 ),
            .clk(N__7110),
            .ce(),
            .sr(N__7001));
    defparam \Instance3.r_Count_16_LC_8_10_7 .C_ON=1'b1;
    defparam \Instance3.r_Count_16_LC_8_10_7 .SEQ_MODE=4'b1000;
    defparam \Instance3.r_Count_16_LC_8_10_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Instance3.r_Count_16_LC_8_10_7  (
            .in0(_gnd_net_),
            .in1(N__7206),
            .in2(_gnd_net_),
            .in3(N__7188),
            .lcout(\Instance3.r_CountZ0Z_16 ),
            .ltout(),
            .carryin(\Instance3.r_Count_2_cry_15 ),
            .carryout(\Instance3.r_Count_2_cry_16 ),
            .clk(N__7110),
            .ce(),
            .sr(N__7001));
    defparam \Instance3.r_Count_17_LC_8_11_0 .C_ON=1'b0;
    defparam \Instance3.r_Count_17_LC_8_11_0 .SEQ_MODE=4'b1000;
    defparam \Instance3.r_Count_17_LC_8_11_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Instance3.r_Count_17_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(N__7182),
            .in2(_gnd_net_),
            .in3(N__7185),
            .lcout(\Instance3.r_CountZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7113),
            .ce(),
            .sr(N__7002));
    defparam \Instance3.r_Count_0_LC_9_10_0 .C_ON=1'b0;
    defparam \Instance3.r_Count_0_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \Instance3.r_Count_0_LC_9_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Instance3.r_Count_0_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7161),
            .lcout(\Instance3.r_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7114),
            .ce(),
            .sr(N__7000));
    defparam \Instance3.r_Count_1_LC_9_10_1 .C_ON=1'b0;
    defparam \Instance3.r_Count_1_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \Instance3.r_Count_1_LC_9_10_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \Instance3.r_Count_1_LC_9_10_1  (
            .in0(N__7162),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7136),
            .lcout(\Instance3.r_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7114),
            .ce(),
            .sr(N__7000));
endmodule // simpleprocessor_top
